module xor_gate (
    input a,
    input b,
    output y
);

 wire net1;
 wire net2;
 wire net3;
 xor2_4 _0_ (.A(net2),
    .B(net1),
    .X(net3));
 decap_3 PHY_EDGE_ROW_0_Right_0 ();
 decap_3 PHY_EDGE_ROW_1_Right_1 ();
 decap_3 PHY_EDGE_ROW_2_Right_2 ();
 decap_3 PHY_EDGE_ROW_3_Right_3 ();
 decap_3 PHY_EDGE_ROW_4_Right_4 ();
 decap_3 PHY_EDGE_ROW_5_Right_5 ();
 decap_3 PHY_EDGE_ROW_6_Right_6 ();
 decap_3 PHY_EDGE_ROW_7_Right_7 ();
 decap_3 PHY_EDGE_ROW_8_Right_8 ();
 decap_3 PHY_EDGE_ROW_9_Right_9 ();
 decap_3 PHY_EDGE_ROW_10_Right_10 ();
 decap_3 PHY_EDGE_ROW_11_Right_11 ();
 decap_3 PHY_EDGE_ROW_12_Right_12 ();
 decap_3 PHY_EDGE_ROW_13_Right_13 ();
 decap_3 PHY_EDGE_ROW_14_Right_14 ();
 decap_3 PHY_EDGE_ROW_15_Right_15 ();
 decap_3 PHY_EDGE_ROW_16_Right_16 ();
 decap_3 PHY_EDGE_ROW_17_Right_17 ();
 decap_3 PHY_EDGE_ROW_18_Right_18 ();
 decap_3 PHY_EDGE_ROW_19_Right_19 ();
 decap_3 PHY_EDGE_ROW_20_Right_20 ();
 decap_3 PHY_EDGE_ROW_21_Right_21 ();
 decap_3 PHY_EDGE_ROW_22_Right_22 ();
 decap_3 PHY_EDGE_ROW_23_Right_23 ();
 decap_3 PHY_EDGE_ROW_24_Right_24 ();
 decap_3 PHY_EDGE_ROW_25_Right_25 ();
 decap_3 PHY_EDGE_ROW_26_Right_26 ();
 decap_3 PHY_EDGE_ROW_27_Right_27 ();
 decap_3 PHY_EDGE_ROW_28_Right_28 ();
 decap_3 PHY_EDGE_ROW_29_Right_29 ();
 decap_3 PHY_EDGE_ROW_30_Right_30 ();
 decap_3 PHY_EDGE_ROW_31_Right_31 ();
 decap_3 PHY_EDGE_ROW_32_Right_32 ();
 decap_3 PHY_EDGE_ROW_33_Right_33 ();
 decap_3 PHY_EDGE_ROW_34_Right_34 ();
 decap_3 PHY_EDGE_ROW_35_Right_35 ();
 decap_3 PHY_EDGE_ROW_36_Right_36 ();
 decap_3 PHY_EDGE_ROW_37_Right_37 ();
 decap_3 PHY_EDGE_ROW_38_Right_38 ();
 decap_3 PHY_EDGE_ROW_39_Right_39 ();
 decap_3 PHY_EDGE_ROW_40_Right_40 ();
 decap_3 PHY_EDGE_ROW_41_Right_41 ();
 decap_3 PHY_EDGE_ROW_42_Right_42 ();
 decap_3 PHY_EDGE_ROW_43_Right_43 ();
 decap_3 PHY_EDGE_ROW_44_Right_44 ();
 decap_3 PHY_EDGE_ROW_45_Right_45 ();
 decap_3 PHY_EDGE_ROW_46_Right_46 ();
 decap_3 PHY_EDGE_ROW_47_Right_47 ();
 decap_3 PHY_EDGE_ROW_48_Right_48 ();
 decap_3 PHY_EDGE_ROW_49_Right_49 ();
 decap_3 PHY_EDGE_ROW_50_Right_50 ();
 decap_3 PHY_EDGE_ROW_51_Right_51 ();
 decap_3 PHY_EDGE_ROW_52_Right_52 ();
 decap_3 PHY_EDGE_ROW_53_Right_53 ();
 decap_3 PHY_EDGE_ROW_54_Right_54 ();
 decap_3 PHY_EDGE_ROW_55_Right_55 ();
 decap_3 PHY_EDGE_ROW_56_Right_56 ();
 decap_3 PHY_EDGE_ROW_57_Right_57 ();
 decap_3 PHY_EDGE_ROW_58_Right_58 ();
 decap_3 PHY_EDGE_ROW_59_Right_59 ();
 decap_3 PHY_EDGE_ROW_60_Right_60 ();
 decap_3 PHY_EDGE_ROW_61_Right_61 ();
 decap_3 PHY_EDGE_ROW_62_Right_62 ();
 decap_3 PHY_EDGE_ROW_63_Right_63 ();
 decap_3 PHY_EDGE_ROW_64_Right_64 ();
 decap_3 PHY_EDGE_ROW_65_Right_65 ();
 decap_3 PHY_EDGE_ROW_66_Right_66 ();
 decap_3 PHY_EDGE_ROW_67_Right_67 ();
 decap_3 PHY_EDGE_ROW_68_Right_68 ();
 decap_3 PHY_EDGE_ROW_69_Right_69 ();
 decap_3 PHY_EDGE_ROW_70_Right_70 ();
 decap_3 PHY_EDGE_ROW_71_Right_71 ();
 decap_3 PHY_EDGE_ROW_72_Right_72 ();
 decap_3 PHY_EDGE_ROW_73_Right_73 ();
 decap_3 PHY_EDGE_ROW_74_Right_74 ();
 decap_3 PHY_EDGE_ROW_75_Right_75 ();
 decap_3 PHY_EDGE_ROW_76_Right_76 ();
 decap_3 PHY_EDGE_ROW_77_Right_77 ();
 decap_3 PHY_EDGE_ROW_78_Right_78 ();
 decap_3 PHY_EDGE_ROW_79_Right_79 ();
 decap_3 PHY_EDGE_ROW_80_Right_80 ();
 decap_3 PHY_EDGE_ROW_81_Right_81 ();
 decap_3 PHY_EDGE_ROW_82_Right_82 ();
 decap_3 PHY_EDGE_ROW_83_Right_83 ();
 decap_3 PHY_EDGE_ROW_84_Right_84 ();
 decap_3 PHY_EDGE_ROW_85_Right_85 ();
 decap_3 PHY_EDGE_ROW_86_Right_86 ();
 decap_3 PHY_EDGE_ROW_87_Right_87 ();
 decap_3 PHY_EDGE_ROW_88_Right_88 ();
 decap_3 PHY_EDGE_ROW_89_Right_89 ();
 decap_3 PHY_EDGE_ROW_90_Right_90 ();
 decap_3 PHY_EDGE_ROW_91_Right_91 ();
 decap_3 PHY_EDGE_ROW_92_Right_92 ();
 decap_3 PHY_EDGE_ROW_93_Right_93 ();
 decap_3 PHY_EDGE_ROW_94_Right_94 ();
 decap_3 PHY_EDGE_ROW_95_Right_95 ();
 decap_3 PHY_EDGE_ROW_96_Right_96 ();
 decap_3 PHY_EDGE_ROW_97_Right_97 ();
 decap_3 PHY_EDGE_ROW_98_Right_98 ();
 decap_3 PHY_EDGE_ROW_99_Right_99 ();
 decap_3 PHY_EDGE_ROW_100_Right_100 ();
 decap_3 PHY_EDGE_ROW_101_Right_101 ();
 decap_3 PHY_EDGE_ROW_0_Left_102 ();
 decap_3 PHY_EDGE_ROW_1_Left_103 ();
 decap_3 PHY_EDGE_ROW_2_Left_104 ();
 decap_3 PHY_EDGE_ROW_3_Left_105 ();
 decap_3 PHY_EDGE_ROW_4_Left_106 ();
 decap_3 PHY_EDGE_ROW_5_Left_107 ();
 decap_3 PHY_EDGE_ROW_6_Left_108 ();
 decap_3 PHY_EDGE_ROW_7_Left_109 ();
 decap_3 PHY_EDGE_ROW_8_Left_110 ();
 decap_3 PHY_EDGE_ROW_9_Left_111 ();
 decap_3 PHY_EDGE_ROW_10_Left_112 ();
 decap_3 PHY_EDGE_ROW_11_Left_113 ();
 decap_3 PHY_EDGE_ROW_12_Left_114 ();
 decap_3 PHY_EDGE_ROW_13_Left_115 ();
 decap_3 PHY_EDGE_ROW_14_Left_116 ();
 decap_3 PHY_EDGE_ROW_15_Left_117 ();
 decap_3 PHY_EDGE_ROW_16_Left_118 ();
 decap_3 PHY_EDGE_ROW_17_Left_119 ();
 decap_3 PHY_EDGE_ROW_18_Left_120 ();
 decap_3 PHY_EDGE_ROW_19_Left_121 ();
 decap_3 PHY_EDGE_ROW_20_Left_122 ();
 decap_3 PHY_EDGE_ROW_21_Left_123 ();
 decap_3 PHY_EDGE_ROW_22_Left_124 ();
 decap_3 PHY_EDGE_ROW_23_Left_125 ();
 decap_3 PHY_EDGE_ROW_24_Left_126 ();
 decap_3 PHY_EDGE_ROW_25_Left_127 ();
 decap_3 PHY_EDGE_ROW_26_Left_128 ();
 decap_3 PHY_EDGE_ROW_27_Left_129 ();
 decap_3 PHY_EDGE_ROW_28_Left_130 ();
 decap_3 PHY_EDGE_ROW_29_Left_131 ();
 decap_3 PHY_EDGE_ROW_30_Left_132 ();
 decap_3 PHY_EDGE_ROW_31_Left_133 ();
 decap_3 PHY_EDGE_ROW_32_Left_134 ();
 decap_3 PHY_EDGE_ROW_33_Left_135 ();
 decap_3 PHY_EDGE_ROW_34_Left_136 ();
 decap_3 PHY_EDGE_ROW_35_Left_137 ();
 decap_3 PHY_EDGE_ROW_36_Left_138 ();
 decap_3 PHY_EDGE_ROW_37_Left_139 ();
 decap_3 PHY_EDGE_ROW_38_Left_140 ();
 decap_3 PHY_EDGE_ROW_39_Left_141 ();
 decap_3 PHY_EDGE_ROW_40_Left_142 ();
 decap_3 PHY_EDGE_ROW_41_Left_143 ();
 decap_3 PHY_EDGE_ROW_42_Left_144 ();
 decap_3 PHY_EDGE_ROW_43_Left_145 ();
 decap_3 PHY_EDGE_ROW_44_Left_146 ();
 decap_3 PHY_EDGE_ROW_45_Left_147 ();
 decap_3 PHY_EDGE_ROW_46_Left_148 ();
 decap_3 PHY_EDGE_ROW_47_Left_149 ();
 decap_3 PHY_EDGE_ROW_48_Left_150 ();
 decap_3 PHY_EDGE_ROW_49_Left_151 ();
 decap_3 PHY_EDGE_ROW_50_Left_152 ();
 decap_3 PHY_EDGE_ROW_51_Left_153 ();
 decap_3 PHY_EDGE_ROW_52_Left_154 ();
 decap_3 PHY_EDGE_ROW_53_Left_155 ();
 decap_3 PHY_EDGE_ROW_54_Left_156 ();
 decap_3 PHY_EDGE_ROW_55_Left_157 ();
 decap_3 PHY_EDGE_ROW_56_Left_158 ();
 decap_3 PHY_EDGE_ROW_57_Left_159 ();
 decap_3 PHY_EDGE_ROW_58_Left_160 ();
 decap_3 PHY_EDGE_ROW_59_Left_161 ();
 decap_3 PHY_EDGE_ROW_60_Left_162 ();
 decap_3 PHY_EDGE_ROW_61_Left_163 ();
 decap_3 PHY_EDGE_ROW_62_Left_164 ();
 decap_3 PHY_EDGE_ROW_63_Left_165 ();
 decap_3 PHY_EDGE_ROW_64_Left_166 ();
 decap_3 PHY_EDGE_ROW_65_Left_167 ();
 decap_3 PHY_EDGE_ROW_66_Left_168 ();
 decap_3 PHY_EDGE_ROW_67_Left_169 ();
 decap_3 PHY_EDGE_ROW_68_Left_170 ();
 decap_3 PHY_EDGE_ROW_69_Left_171 ();
 decap_3 PHY_EDGE_ROW_70_Left_172 ();
 decap_3 PHY_EDGE_ROW_71_Left_173 ();
 decap_3 PHY_EDGE_ROW_72_Left_174 ();
 decap_3 PHY_EDGE_ROW_73_Left_175 ();
 decap_3 PHY_EDGE_ROW_74_Left_176 ();
 decap_3 PHY_EDGE_ROW_75_Left_177 ();
 decap_3 PHY_EDGE_ROW_76_Left_178 ();
 decap_3 PHY_EDGE_ROW_77_Left_179 ();
 decap_3 PHY_EDGE_ROW_78_Left_180 ();
 decap_3 PHY_EDGE_ROW_79_Left_181 ();
 decap_3 PHY_EDGE_ROW_80_Left_182 ();
 decap_3 PHY_EDGE_ROW_81_Left_183 ();
 decap_3 PHY_EDGE_ROW_82_Left_184 ();
 decap_3 PHY_EDGE_ROW_83_Left_185 ();
 decap_3 PHY_EDGE_ROW_84_Left_186 ();
 decap_3 PHY_EDGE_ROW_85_Left_187 ();
 decap_3 PHY_EDGE_ROW_86_Left_188 ();
 decap_3 PHY_EDGE_ROW_87_Left_189 ();
 decap_3 PHY_EDGE_ROW_88_Left_190 ();
 decap_3 PHY_EDGE_ROW_89_Left_191 ();
 decap_3 PHY_EDGE_ROW_90_Left_192 ();
 decap_3 PHY_EDGE_ROW_91_Left_193 ();
 decap_3 PHY_EDGE_ROW_92_Left_194 ();
 decap_3 PHY_EDGE_ROW_93_Left_195 ();
 decap_3 PHY_EDGE_ROW_94_Left_196 ();
 decap_3 PHY_EDGE_ROW_95_Left_197 ();
 decap_3 PHY_EDGE_ROW_96_Left_198 ();
 decap_3 PHY_EDGE_ROW_97_Left_199 ();
 decap_3 PHY_EDGE_ROW_98_Left_200 ();
 decap_3 PHY_EDGE_ROW_99_Left_201 ();
 decap_3 PHY_EDGE_ROW_100_Left_202 ();
 decap_3 PHY_EDGE_ROW_101_Left_203 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 dlymetal6s2s_1 input1 (.A(a),
    .X(net1));
 clkbuf_2 input2 (.A(b),
    .X(net2));
 buf_2 output3 (.A(net3),
    .X(y));
 decap_12 FILLER_0_3 ();
 decap_12 FILLER_0_15 ();
 fill_1 FILLER_0_27 ();
 decap_12 FILLER_0_29 ();
 decap_12 FILLER_0_41 ();
 fill_2 FILLER_0_53 ();
 fill_1 FILLER_0_55 ();
 decap_12 FILLER_0_57 ();
 decap_12 FILLER_0_69 ();
 fill_2 FILLER_0_81 ();
 fill_1 FILLER_0_83 ();
 decap_12 FILLER_0_85 ();
 decap_12 FILLER_0_97 ();
 fill_2 FILLER_0_109 ();
 fill_1 FILLER_0_111 ();
 decap_12 FILLER_0_113 ();
 decap_12 FILLER_0_125 ();
 fill_2 FILLER_0_137 ();
 fill_1 FILLER_0_139 ();
 decap_12 FILLER_0_141 ();
 decap_12 FILLER_0_153 ();
 fill_2 FILLER_0_165 ();
 fill_1 FILLER_0_167 ();
 decap_12 FILLER_0_169 ();
 decap_12 FILLER_0_181 ();
 fill_2 FILLER_0_193 ();
 fill_1 FILLER_0_195 ();
 decap_12 FILLER_0_197 ();
 decap_12 FILLER_0_209 ();
 fill_2 FILLER_0_221 ();
 fill_1 FILLER_0_223 ();
 decap_12 FILLER_0_225 ();
 decap_12 FILLER_0_237 ();
 fill_2 FILLER_0_249 ();
 fill_1 FILLER_0_251 ();
 decap_12 FILLER_0_253 ();
 decap_12 FILLER_0_265 ();
 fill_2 FILLER_0_277 ();
 fill_1 FILLER_0_279 ();
 decap_12 FILLER_0_281 ();
 decap_12 FILLER_0_293 ();
 fill_2 FILLER_0_305 ();
 fill_1 FILLER_0_307 ();
 decap_12 FILLER_0_309 ();
 decap_12 FILLER_0_321 ();
 fill_2 FILLER_0_333 ();
 fill_1 FILLER_0_335 ();
 decap_12 FILLER_0_337 ();
 decap_12 FILLER_0_349 ();
 fill_2 FILLER_0_361 ();
 fill_1 FILLER_0_363 ();
 decap_12 FILLER_0_365 ();
 decap_12 FILLER_0_377 ();
 fill_2 FILLER_0_389 ();
 fill_1 FILLER_0_391 ();
 decap_12 FILLER_0_393 ();
 decap_12 FILLER_0_405 ();
 fill_2 FILLER_0_417 ();
 fill_1 FILLER_0_419 ();
 decap_12 FILLER_0_421 ();
 decap_12 FILLER_0_433 ();
 fill_2 FILLER_0_445 ();
 fill_1 FILLER_0_447 ();
 decap_12 FILLER_0_449 ();
 decap_12 FILLER_0_461 ();
 fill_2 FILLER_0_473 ();
 fill_1 FILLER_0_475 ();
 decap_12 FILLER_0_477 ();
 decap_12 FILLER_0_489 ();
 fill_2 FILLER_0_501 ();
 fill_1 FILLER_0_503 ();
 decap_12 FILLER_0_505 ();
 decap_12 FILLER_0_517 ();
 fill_2 FILLER_0_529 ();
 fill_1 FILLER_0_531 ();
 decap_12 FILLER_0_533 ();
 decap_12 FILLER_0_545 ();
 fill_2 FILLER_0_557 ();
 fill_1 FILLER_0_559 ();
 decap_12 FILLER_0_561 ();
 decap_12 FILLER_0_573 ();
 fill_2 FILLER_0_585 ();
 fill_1 FILLER_0_587 ();
 decap_12 FILLER_0_589 ();
 decap_12 FILLER_0_601 ();
 fill_2 FILLER_0_613 ();
 fill_1 FILLER_0_615 ();
 fill_8 FILLER_0_617 ();
 decap_12 FILLER_1_3 ();
 decap_12 FILLER_1_15 ();
 decap_12 FILLER_1_27 ();
 decap_12 FILLER_1_39 ();
 fill_4 FILLER_1_51 ();
 fill_1 FILLER_1_55 ();
 decap_12 FILLER_1_57 ();
 decap_12 FILLER_1_69 ();
 decap_12 FILLER_1_81 ();
 decap_12 FILLER_1_93 ();
 fill_4 FILLER_1_105 ();
 fill_2 FILLER_1_109 ();
 fill_1 FILLER_1_111 ();
 decap_12 FILLER_1_113 ();
 decap_12 FILLER_1_125 ();
 decap_12 FILLER_1_137 ();
 decap_12 FILLER_1_149 ();
 fill_4 FILLER_1_161 ();
 fill_2 FILLER_1_165 ();
 fill_1 FILLER_1_167 ();
 decap_12 FILLER_1_169 ();
 decap_12 FILLER_1_181 ();
 decap_12 FILLER_1_193 ();
 decap_12 FILLER_1_205 ();
 fill_4 FILLER_1_217 ();
 fill_2 FILLER_1_221 ();
 fill_1 FILLER_1_223 ();
 decap_12 FILLER_1_225 ();
 decap_12 FILLER_1_237 ();
 decap_12 FILLER_1_249 ();
 decap_12 FILLER_1_261 ();
 fill_4 FILLER_1_273 ();
 fill_2 FILLER_1_277 ();
 fill_1 FILLER_1_279 ();
 decap_12 FILLER_1_281 ();
 decap_12 FILLER_1_293 ();
 decap_12 FILLER_1_305 ();
 decap_12 FILLER_1_317 ();
 fill_4 FILLER_1_329 ();
 fill_2 FILLER_1_333 ();
 fill_1 FILLER_1_335 ();
 decap_12 FILLER_1_337 ();
 decap_12 FILLER_1_349 ();
 decap_12 FILLER_1_361 ();
 decap_12 FILLER_1_373 ();
 fill_4 FILLER_1_385 ();
 fill_2 FILLER_1_389 ();
 fill_1 FILLER_1_391 ();
 decap_12 FILLER_1_393 ();
 decap_12 FILLER_1_405 ();
 decap_12 FILLER_1_417 ();
 decap_12 FILLER_1_429 ();
 fill_4 FILLER_1_441 ();
 fill_2 FILLER_1_445 ();
 fill_1 FILLER_1_447 ();
 decap_12 FILLER_1_449 ();
 decap_12 FILLER_1_461 ();
 decap_12 FILLER_1_473 ();
 decap_12 FILLER_1_485 ();
 fill_4 FILLER_1_497 ();
 fill_2 FILLER_1_501 ();
 fill_1 FILLER_1_503 ();
 decap_12 FILLER_1_505 ();
 decap_12 FILLER_1_517 ();
 decap_12 FILLER_1_529 ();
 decap_12 FILLER_1_541 ();
 fill_4 FILLER_1_553 ();
 fill_2 FILLER_1_557 ();
 fill_1 FILLER_1_559 ();
 decap_12 FILLER_1_561 ();
 decap_12 FILLER_1_573 ();
 decap_12 FILLER_1_585 ();
 decap_12 FILLER_1_597 ();
 fill_4 FILLER_1_609 ();
 fill_2 FILLER_1_613 ();
 fill_1 FILLER_1_615 ();
 fill_8 FILLER_1_617 ();
 decap_12 FILLER_2_3 ();
 decap_12 FILLER_2_15 ();
 fill_1 FILLER_2_27 ();
 decap_12 FILLER_2_29 ();
 decap_12 FILLER_2_41 ();
 decap_12 FILLER_2_53 ();
 decap_12 FILLER_2_65 ();
 fill_4 FILLER_2_77 ();
 fill_2 FILLER_2_81 ();
 fill_1 FILLER_2_83 ();
 decap_12 FILLER_2_85 ();
 decap_12 FILLER_2_97 ();
 decap_12 FILLER_2_109 ();
 decap_12 FILLER_2_121 ();
 fill_4 FILLER_2_133 ();
 fill_2 FILLER_2_137 ();
 fill_1 FILLER_2_139 ();
 decap_12 FILLER_2_141 ();
 decap_12 FILLER_2_153 ();
 decap_12 FILLER_2_165 ();
 decap_12 FILLER_2_177 ();
 fill_4 FILLER_2_189 ();
 fill_2 FILLER_2_193 ();
 fill_1 FILLER_2_195 ();
 decap_12 FILLER_2_197 ();
 decap_12 FILLER_2_209 ();
 decap_12 FILLER_2_221 ();
 decap_12 FILLER_2_233 ();
 fill_4 FILLER_2_245 ();
 fill_2 FILLER_2_249 ();
 fill_1 FILLER_2_251 ();
 decap_12 FILLER_2_253 ();
 decap_12 FILLER_2_265 ();
 decap_12 FILLER_2_277 ();
 decap_12 FILLER_2_289 ();
 fill_4 FILLER_2_301 ();
 fill_2 FILLER_2_305 ();
 fill_1 FILLER_2_307 ();
 decap_12 FILLER_2_309 ();
 decap_12 FILLER_2_321 ();
 decap_12 FILLER_2_333 ();
 decap_12 FILLER_2_345 ();
 fill_4 FILLER_2_357 ();
 fill_2 FILLER_2_361 ();
 fill_1 FILLER_2_363 ();
 decap_12 FILLER_2_365 ();
 decap_12 FILLER_2_377 ();
 decap_12 FILLER_2_389 ();
 decap_12 FILLER_2_401 ();
 fill_4 FILLER_2_413 ();
 fill_2 FILLER_2_417 ();
 fill_1 FILLER_2_419 ();
 decap_12 FILLER_2_421 ();
 decap_12 FILLER_2_433 ();
 decap_12 FILLER_2_445 ();
 decap_12 FILLER_2_457 ();
 fill_4 FILLER_2_469 ();
 fill_2 FILLER_2_473 ();
 fill_1 FILLER_2_475 ();
 decap_12 FILLER_2_477 ();
 decap_12 FILLER_2_489 ();
 decap_12 FILLER_2_501 ();
 decap_12 FILLER_2_513 ();
 fill_4 FILLER_2_525 ();
 fill_2 FILLER_2_529 ();
 fill_1 FILLER_2_531 ();
 decap_12 FILLER_2_533 ();
 decap_12 FILLER_2_545 ();
 decap_12 FILLER_2_557 ();
 decap_12 FILLER_2_569 ();
 fill_4 FILLER_2_581 ();
 fill_2 FILLER_2_585 ();
 fill_1 FILLER_2_587 ();
 decap_12 FILLER_2_589 ();
 decap_12 FILLER_2_601 ();
 decap_12 FILLER_2_613 ();
 decap_12 FILLER_3_3 ();
 decap_12 FILLER_3_15 ();
 decap_12 FILLER_3_27 ();
 decap_12 FILLER_3_39 ();
 fill_4 FILLER_3_51 ();
 fill_1 FILLER_3_55 ();
 decap_12 FILLER_3_57 ();
 decap_12 FILLER_3_69 ();
 decap_12 FILLER_3_81 ();
 decap_12 FILLER_3_93 ();
 fill_4 FILLER_3_105 ();
 fill_2 FILLER_3_109 ();
 fill_1 FILLER_3_111 ();
 decap_12 FILLER_3_113 ();
 decap_12 FILLER_3_125 ();
 decap_12 FILLER_3_137 ();
 decap_12 FILLER_3_149 ();
 fill_4 FILLER_3_161 ();
 fill_2 FILLER_3_165 ();
 fill_1 FILLER_3_167 ();
 decap_12 FILLER_3_169 ();
 decap_12 FILLER_3_181 ();
 decap_12 FILLER_3_193 ();
 decap_12 FILLER_3_205 ();
 fill_4 FILLER_3_217 ();
 fill_2 FILLER_3_221 ();
 fill_1 FILLER_3_223 ();
 decap_12 FILLER_3_225 ();
 decap_12 FILLER_3_237 ();
 decap_12 FILLER_3_249 ();
 decap_12 FILLER_3_261 ();
 fill_4 FILLER_3_273 ();
 fill_2 FILLER_3_277 ();
 fill_1 FILLER_3_279 ();
 decap_12 FILLER_3_281 ();
 decap_12 FILLER_3_293 ();
 decap_12 FILLER_3_305 ();
 decap_12 FILLER_3_317 ();
 fill_4 FILLER_3_329 ();
 fill_2 FILLER_3_333 ();
 fill_1 FILLER_3_335 ();
 decap_12 FILLER_3_337 ();
 decap_12 FILLER_3_349 ();
 decap_12 FILLER_3_361 ();
 decap_12 FILLER_3_373 ();
 fill_4 FILLER_3_385 ();
 fill_2 FILLER_3_389 ();
 fill_1 FILLER_3_391 ();
 decap_12 FILLER_3_393 ();
 decap_12 FILLER_3_405 ();
 decap_12 FILLER_3_417 ();
 decap_12 FILLER_3_429 ();
 fill_4 FILLER_3_441 ();
 fill_2 FILLER_3_445 ();
 fill_1 FILLER_3_447 ();
 decap_12 FILLER_3_449 ();
 decap_12 FILLER_3_461 ();
 decap_12 FILLER_3_473 ();
 decap_12 FILLER_3_485 ();
 fill_4 FILLER_3_497 ();
 fill_2 FILLER_3_501 ();
 fill_1 FILLER_3_503 ();
 decap_12 FILLER_3_505 ();
 decap_12 FILLER_3_517 ();
 decap_12 FILLER_3_529 ();
 decap_12 FILLER_3_541 ();
 fill_4 FILLER_3_553 ();
 fill_2 FILLER_3_557 ();
 fill_1 FILLER_3_559 ();
 decap_12 FILLER_3_561 ();
 decap_12 FILLER_3_573 ();
 decap_12 FILLER_3_585 ();
 decap_12 FILLER_3_597 ();
 fill_4 FILLER_3_609 ();
 fill_2 FILLER_3_613 ();
 fill_1 FILLER_3_615 ();
 fill_8 FILLER_3_617 ();
 decap_12 FILLER_4_3 ();
 decap_12 FILLER_4_15 ();
 fill_1 FILLER_4_27 ();
 decap_12 FILLER_4_29 ();
 decap_12 FILLER_4_41 ();
 decap_12 FILLER_4_53 ();
 decap_12 FILLER_4_65 ();
 fill_4 FILLER_4_77 ();
 fill_2 FILLER_4_81 ();
 fill_1 FILLER_4_83 ();
 decap_12 FILLER_4_85 ();
 decap_12 FILLER_4_97 ();
 decap_12 FILLER_4_109 ();
 decap_12 FILLER_4_121 ();
 fill_4 FILLER_4_133 ();
 fill_2 FILLER_4_137 ();
 fill_1 FILLER_4_139 ();
 decap_12 FILLER_4_141 ();
 decap_12 FILLER_4_153 ();
 decap_12 FILLER_4_165 ();
 decap_12 FILLER_4_177 ();
 fill_4 FILLER_4_189 ();
 fill_2 FILLER_4_193 ();
 fill_1 FILLER_4_195 ();
 decap_12 FILLER_4_197 ();
 decap_12 FILLER_4_209 ();
 decap_12 FILLER_4_221 ();
 decap_12 FILLER_4_233 ();
 fill_4 FILLER_4_245 ();
 fill_2 FILLER_4_249 ();
 fill_1 FILLER_4_251 ();
 decap_12 FILLER_4_253 ();
 decap_12 FILLER_4_265 ();
 decap_12 FILLER_4_277 ();
 decap_12 FILLER_4_289 ();
 fill_4 FILLER_4_301 ();
 fill_2 FILLER_4_305 ();
 fill_1 FILLER_4_307 ();
 decap_12 FILLER_4_309 ();
 decap_12 FILLER_4_321 ();
 decap_12 FILLER_4_333 ();
 decap_12 FILLER_4_345 ();
 fill_4 FILLER_4_357 ();
 fill_2 FILLER_4_361 ();
 fill_1 FILLER_4_363 ();
 decap_12 FILLER_4_365 ();
 decap_12 FILLER_4_377 ();
 decap_12 FILLER_4_389 ();
 decap_12 FILLER_4_401 ();
 fill_4 FILLER_4_413 ();
 fill_2 FILLER_4_417 ();
 fill_1 FILLER_4_419 ();
 decap_12 FILLER_4_421 ();
 decap_12 FILLER_4_433 ();
 decap_12 FILLER_4_445 ();
 decap_12 FILLER_4_457 ();
 fill_4 FILLER_4_469 ();
 fill_2 FILLER_4_473 ();
 fill_1 FILLER_4_475 ();
 decap_12 FILLER_4_477 ();
 decap_12 FILLER_4_489 ();
 decap_12 FILLER_4_501 ();
 decap_12 FILLER_4_513 ();
 fill_4 FILLER_4_525 ();
 fill_2 FILLER_4_529 ();
 fill_1 FILLER_4_531 ();
 decap_12 FILLER_4_533 ();
 decap_12 FILLER_4_545 ();
 decap_12 FILLER_4_557 ();
 decap_12 FILLER_4_569 ();
 fill_4 FILLER_4_581 ();
 fill_2 FILLER_4_585 ();
 fill_1 FILLER_4_587 ();
 decap_12 FILLER_4_589 ();
 decap_12 FILLER_4_601 ();
 decap_12 FILLER_4_613 ();
 decap_12 FILLER_5_3 ();
 decap_12 FILLER_5_15 ();
 decap_12 FILLER_5_27 ();
 decap_12 FILLER_5_39 ();
 fill_4 FILLER_5_51 ();
 fill_1 FILLER_5_55 ();
 decap_12 FILLER_5_57 ();
 decap_12 FILLER_5_69 ();
 decap_12 FILLER_5_81 ();
 decap_12 FILLER_5_93 ();
 fill_4 FILLER_5_105 ();
 fill_2 FILLER_5_109 ();
 fill_1 FILLER_5_111 ();
 decap_12 FILLER_5_113 ();
 decap_12 FILLER_5_125 ();
 decap_12 FILLER_5_137 ();
 decap_12 FILLER_5_149 ();
 fill_4 FILLER_5_161 ();
 fill_2 FILLER_5_165 ();
 fill_1 FILLER_5_167 ();
 decap_12 FILLER_5_169 ();
 decap_12 FILLER_5_181 ();
 decap_12 FILLER_5_193 ();
 decap_12 FILLER_5_205 ();
 fill_4 FILLER_5_217 ();
 fill_2 FILLER_5_221 ();
 fill_1 FILLER_5_223 ();
 decap_12 FILLER_5_225 ();
 decap_12 FILLER_5_237 ();
 decap_12 FILLER_5_249 ();
 decap_12 FILLER_5_261 ();
 fill_4 FILLER_5_273 ();
 fill_2 FILLER_5_277 ();
 fill_1 FILLER_5_279 ();
 decap_12 FILLER_5_281 ();
 decap_12 FILLER_5_293 ();
 decap_12 FILLER_5_305 ();
 decap_12 FILLER_5_317 ();
 fill_4 FILLER_5_329 ();
 fill_2 FILLER_5_333 ();
 fill_1 FILLER_5_335 ();
 decap_12 FILLER_5_337 ();
 decap_12 FILLER_5_349 ();
 decap_12 FILLER_5_361 ();
 decap_12 FILLER_5_373 ();
 fill_4 FILLER_5_385 ();
 fill_2 FILLER_5_389 ();
 fill_1 FILLER_5_391 ();
 decap_12 FILLER_5_393 ();
 decap_12 FILLER_5_405 ();
 decap_12 FILLER_5_417 ();
 decap_12 FILLER_5_429 ();
 fill_4 FILLER_5_441 ();
 fill_2 FILLER_5_445 ();
 fill_1 FILLER_5_447 ();
 decap_12 FILLER_5_449 ();
 decap_12 FILLER_5_461 ();
 decap_12 FILLER_5_473 ();
 decap_12 FILLER_5_485 ();
 fill_4 FILLER_5_497 ();
 fill_2 FILLER_5_501 ();
 fill_1 FILLER_5_503 ();
 decap_12 FILLER_5_505 ();
 decap_12 FILLER_5_517 ();
 decap_12 FILLER_5_529 ();
 decap_12 FILLER_5_541 ();
 fill_4 FILLER_5_553 ();
 fill_2 FILLER_5_557 ();
 fill_1 FILLER_5_559 ();
 decap_12 FILLER_5_561 ();
 decap_12 FILLER_5_573 ();
 decap_12 FILLER_5_585 ();
 decap_12 FILLER_5_597 ();
 fill_4 FILLER_5_609 ();
 fill_2 FILLER_5_613 ();
 fill_1 FILLER_5_615 ();
 fill_8 FILLER_5_617 ();
 decap_12 FILLER_6_3 ();
 decap_12 FILLER_6_15 ();
 fill_1 FILLER_6_27 ();
 decap_12 FILLER_6_29 ();
 decap_12 FILLER_6_41 ();
 decap_12 FILLER_6_53 ();
 decap_12 FILLER_6_65 ();
 fill_4 FILLER_6_77 ();
 fill_2 FILLER_6_81 ();
 fill_1 FILLER_6_83 ();
 decap_12 FILLER_6_85 ();
 decap_12 FILLER_6_97 ();
 decap_12 FILLER_6_109 ();
 decap_12 FILLER_6_121 ();
 fill_4 FILLER_6_133 ();
 fill_2 FILLER_6_137 ();
 fill_1 FILLER_6_139 ();
 decap_12 FILLER_6_141 ();
 decap_12 FILLER_6_153 ();
 decap_12 FILLER_6_165 ();
 decap_12 FILLER_6_177 ();
 fill_4 FILLER_6_189 ();
 fill_2 FILLER_6_193 ();
 fill_1 FILLER_6_195 ();
 decap_12 FILLER_6_197 ();
 decap_12 FILLER_6_209 ();
 decap_12 FILLER_6_221 ();
 decap_12 FILLER_6_233 ();
 fill_4 FILLER_6_245 ();
 fill_2 FILLER_6_249 ();
 fill_1 FILLER_6_251 ();
 decap_12 FILLER_6_253 ();
 decap_12 FILLER_6_265 ();
 decap_12 FILLER_6_277 ();
 decap_12 FILLER_6_289 ();
 fill_4 FILLER_6_301 ();
 fill_2 FILLER_6_305 ();
 fill_1 FILLER_6_307 ();
 decap_12 FILLER_6_309 ();
 decap_12 FILLER_6_321 ();
 decap_12 FILLER_6_333 ();
 decap_12 FILLER_6_345 ();
 fill_4 FILLER_6_357 ();
 fill_2 FILLER_6_361 ();
 fill_1 FILLER_6_363 ();
 decap_12 FILLER_6_365 ();
 decap_12 FILLER_6_377 ();
 decap_12 FILLER_6_389 ();
 decap_12 FILLER_6_401 ();
 fill_4 FILLER_6_413 ();
 fill_2 FILLER_6_417 ();
 fill_1 FILLER_6_419 ();
 decap_12 FILLER_6_421 ();
 decap_12 FILLER_6_433 ();
 decap_12 FILLER_6_445 ();
 decap_12 FILLER_6_457 ();
 fill_4 FILLER_6_469 ();
 fill_2 FILLER_6_473 ();
 fill_1 FILLER_6_475 ();
 decap_12 FILLER_6_477 ();
 decap_12 FILLER_6_489 ();
 decap_12 FILLER_6_501 ();
 decap_12 FILLER_6_513 ();
 fill_4 FILLER_6_525 ();
 fill_2 FILLER_6_529 ();
 fill_1 FILLER_6_531 ();
 decap_12 FILLER_6_533 ();
 decap_12 FILLER_6_545 ();
 decap_12 FILLER_6_557 ();
 decap_12 FILLER_6_569 ();
 fill_4 FILLER_6_581 ();
 fill_2 FILLER_6_585 ();
 fill_1 FILLER_6_587 ();
 decap_12 FILLER_6_589 ();
 decap_12 FILLER_6_601 ();
 decap_12 FILLER_6_613 ();
 decap_12 FILLER_7_3 ();
 decap_12 FILLER_7_15 ();
 decap_12 FILLER_7_27 ();
 decap_12 FILLER_7_39 ();
 fill_4 FILLER_7_51 ();
 fill_1 FILLER_7_55 ();
 decap_12 FILLER_7_57 ();
 decap_12 FILLER_7_69 ();
 decap_12 FILLER_7_81 ();
 decap_12 FILLER_7_93 ();
 fill_4 FILLER_7_105 ();
 fill_2 FILLER_7_109 ();
 fill_1 FILLER_7_111 ();
 decap_12 FILLER_7_113 ();
 decap_12 FILLER_7_125 ();
 decap_12 FILLER_7_137 ();
 decap_12 FILLER_7_149 ();
 fill_4 FILLER_7_161 ();
 fill_2 FILLER_7_165 ();
 fill_1 FILLER_7_167 ();
 decap_12 FILLER_7_169 ();
 decap_12 FILLER_7_181 ();
 decap_12 FILLER_7_193 ();
 decap_12 FILLER_7_205 ();
 fill_4 FILLER_7_217 ();
 fill_2 FILLER_7_221 ();
 fill_1 FILLER_7_223 ();
 decap_12 FILLER_7_225 ();
 decap_12 FILLER_7_237 ();
 decap_12 FILLER_7_249 ();
 decap_12 FILLER_7_261 ();
 fill_4 FILLER_7_273 ();
 fill_2 FILLER_7_277 ();
 fill_1 FILLER_7_279 ();
 decap_12 FILLER_7_281 ();
 decap_12 FILLER_7_293 ();
 decap_12 FILLER_7_305 ();
 decap_12 FILLER_7_317 ();
 fill_4 FILLER_7_329 ();
 fill_2 FILLER_7_333 ();
 fill_1 FILLER_7_335 ();
 decap_12 FILLER_7_337 ();
 decap_12 FILLER_7_349 ();
 decap_12 FILLER_7_361 ();
 decap_12 FILLER_7_373 ();
 fill_4 FILLER_7_385 ();
 fill_2 FILLER_7_389 ();
 fill_1 FILLER_7_391 ();
 decap_12 FILLER_7_393 ();
 decap_12 FILLER_7_405 ();
 decap_12 FILLER_7_417 ();
 decap_12 FILLER_7_429 ();
 fill_4 FILLER_7_441 ();
 fill_2 FILLER_7_445 ();
 fill_1 FILLER_7_447 ();
 decap_12 FILLER_7_449 ();
 decap_12 FILLER_7_461 ();
 decap_12 FILLER_7_473 ();
 decap_12 FILLER_7_485 ();
 fill_4 FILLER_7_497 ();
 fill_2 FILLER_7_501 ();
 fill_1 FILLER_7_503 ();
 decap_12 FILLER_7_505 ();
 decap_12 FILLER_7_517 ();
 decap_12 FILLER_7_529 ();
 decap_12 FILLER_7_541 ();
 fill_4 FILLER_7_553 ();
 fill_2 FILLER_7_557 ();
 fill_1 FILLER_7_559 ();
 decap_12 FILLER_7_561 ();
 decap_12 FILLER_7_573 ();
 decap_12 FILLER_7_585 ();
 decap_12 FILLER_7_597 ();
 fill_4 FILLER_7_609 ();
 fill_2 FILLER_7_613 ();
 fill_1 FILLER_7_615 ();
 fill_8 FILLER_7_617 ();
 decap_12 FILLER_8_3 ();
 decap_12 FILLER_8_15 ();
 fill_1 FILLER_8_27 ();
 decap_12 FILLER_8_29 ();
 decap_12 FILLER_8_41 ();
 decap_12 FILLER_8_53 ();
 decap_12 FILLER_8_65 ();
 fill_4 FILLER_8_77 ();
 fill_2 FILLER_8_81 ();
 fill_1 FILLER_8_83 ();
 decap_12 FILLER_8_85 ();
 decap_12 FILLER_8_97 ();
 decap_12 FILLER_8_109 ();
 decap_12 FILLER_8_121 ();
 fill_4 FILLER_8_133 ();
 fill_2 FILLER_8_137 ();
 fill_1 FILLER_8_139 ();
 decap_12 FILLER_8_141 ();
 decap_12 FILLER_8_153 ();
 decap_12 FILLER_8_165 ();
 decap_12 FILLER_8_177 ();
 fill_4 FILLER_8_189 ();
 fill_2 FILLER_8_193 ();
 fill_1 FILLER_8_195 ();
 decap_12 FILLER_8_197 ();
 decap_12 FILLER_8_209 ();
 decap_12 FILLER_8_221 ();
 decap_12 FILLER_8_233 ();
 fill_4 FILLER_8_245 ();
 fill_2 FILLER_8_249 ();
 fill_1 FILLER_8_251 ();
 decap_12 FILLER_8_253 ();
 decap_12 FILLER_8_265 ();
 decap_12 FILLER_8_277 ();
 decap_12 FILLER_8_289 ();
 fill_4 FILLER_8_301 ();
 fill_2 FILLER_8_305 ();
 fill_1 FILLER_8_307 ();
 decap_12 FILLER_8_309 ();
 decap_12 FILLER_8_321 ();
 decap_12 FILLER_8_333 ();
 decap_12 FILLER_8_345 ();
 fill_4 FILLER_8_357 ();
 fill_2 FILLER_8_361 ();
 fill_1 FILLER_8_363 ();
 decap_12 FILLER_8_365 ();
 decap_12 FILLER_8_377 ();
 decap_12 FILLER_8_389 ();
 decap_12 FILLER_8_401 ();
 fill_4 FILLER_8_413 ();
 fill_2 FILLER_8_417 ();
 fill_1 FILLER_8_419 ();
 decap_12 FILLER_8_421 ();
 decap_12 FILLER_8_433 ();
 decap_12 FILLER_8_445 ();
 decap_12 FILLER_8_457 ();
 fill_4 FILLER_8_469 ();
 fill_2 FILLER_8_473 ();
 fill_1 FILLER_8_475 ();
 decap_12 FILLER_8_477 ();
 decap_12 FILLER_8_489 ();
 decap_12 FILLER_8_501 ();
 decap_12 FILLER_8_513 ();
 fill_4 FILLER_8_525 ();
 fill_2 FILLER_8_529 ();
 fill_1 FILLER_8_531 ();
 decap_12 FILLER_8_533 ();
 decap_12 FILLER_8_545 ();
 decap_12 FILLER_8_557 ();
 decap_12 FILLER_8_569 ();
 fill_4 FILLER_8_581 ();
 fill_2 FILLER_8_585 ();
 fill_1 FILLER_8_587 ();
 decap_12 FILLER_8_589 ();
 decap_12 FILLER_8_601 ();
 decap_12 FILLER_8_613 ();
 decap_12 FILLER_9_3 ();
 decap_12 FILLER_9_15 ();
 decap_12 FILLER_9_27 ();
 decap_12 FILLER_9_39 ();
 fill_4 FILLER_9_51 ();
 fill_1 FILLER_9_55 ();
 decap_12 FILLER_9_57 ();
 decap_12 FILLER_9_69 ();
 decap_12 FILLER_9_81 ();
 decap_12 FILLER_9_93 ();
 fill_4 FILLER_9_105 ();
 fill_2 FILLER_9_109 ();
 fill_1 FILLER_9_111 ();
 decap_12 FILLER_9_113 ();
 decap_12 FILLER_9_125 ();
 decap_12 FILLER_9_137 ();
 decap_12 FILLER_9_149 ();
 fill_4 FILLER_9_161 ();
 fill_2 FILLER_9_165 ();
 fill_1 FILLER_9_167 ();
 decap_12 FILLER_9_169 ();
 decap_12 FILLER_9_181 ();
 decap_12 FILLER_9_193 ();
 decap_12 FILLER_9_205 ();
 fill_4 FILLER_9_217 ();
 fill_2 FILLER_9_221 ();
 fill_1 FILLER_9_223 ();
 decap_12 FILLER_9_225 ();
 decap_12 FILLER_9_237 ();
 decap_12 FILLER_9_249 ();
 decap_12 FILLER_9_261 ();
 fill_4 FILLER_9_273 ();
 fill_2 FILLER_9_277 ();
 fill_1 FILLER_9_279 ();
 decap_12 FILLER_9_281 ();
 decap_12 FILLER_9_293 ();
 decap_12 FILLER_9_305 ();
 decap_12 FILLER_9_317 ();
 fill_4 FILLER_9_329 ();
 fill_2 FILLER_9_333 ();
 fill_1 FILLER_9_335 ();
 decap_12 FILLER_9_337 ();
 decap_12 FILLER_9_349 ();
 decap_12 FILLER_9_361 ();
 decap_12 FILLER_9_373 ();
 fill_4 FILLER_9_385 ();
 fill_2 FILLER_9_389 ();
 fill_1 FILLER_9_391 ();
 decap_12 FILLER_9_393 ();
 decap_12 FILLER_9_405 ();
 decap_12 FILLER_9_417 ();
 decap_12 FILLER_9_429 ();
 fill_4 FILLER_9_441 ();
 fill_2 FILLER_9_445 ();
 fill_1 FILLER_9_447 ();
 decap_12 FILLER_9_449 ();
 decap_12 FILLER_9_461 ();
 decap_12 FILLER_9_473 ();
 decap_12 FILLER_9_485 ();
 fill_4 FILLER_9_497 ();
 fill_2 FILLER_9_501 ();
 fill_1 FILLER_9_503 ();
 decap_12 FILLER_9_505 ();
 decap_12 FILLER_9_517 ();
 decap_12 FILLER_9_529 ();
 decap_12 FILLER_9_541 ();
 fill_4 FILLER_9_553 ();
 fill_2 FILLER_9_557 ();
 fill_1 FILLER_9_559 ();
 decap_12 FILLER_9_561 ();
 decap_12 FILLER_9_573 ();
 decap_12 FILLER_9_585 ();
 decap_12 FILLER_9_597 ();
 fill_4 FILLER_9_609 ();
 fill_2 FILLER_9_613 ();
 fill_1 FILLER_9_615 ();
 fill_8 FILLER_9_617 ();
 decap_12 FILLER_10_3 ();
 decap_12 FILLER_10_15 ();
 fill_1 FILLER_10_27 ();
 decap_12 FILLER_10_29 ();
 decap_12 FILLER_10_41 ();
 decap_12 FILLER_10_53 ();
 decap_12 FILLER_10_65 ();
 fill_4 FILLER_10_77 ();
 fill_2 FILLER_10_81 ();
 fill_1 FILLER_10_83 ();
 decap_12 FILLER_10_85 ();
 decap_12 FILLER_10_97 ();
 decap_12 FILLER_10_109 ();
 decap_12 FILLER_10_121 ();
 fill_4 FILLER_10_133 ();
 fill_2 FILLER_10_137 ();
 fill_1 FILLER_10_139 ();
 decap_12 FILLER_10_141 ();
 decap_12 FILLER_10_153 ();
 decap_12 FILLER_10_165 ();
 decap_12 FILLER_10_177 ();
 fill_4 FILLER_10_189 ();
 fill_2 FILLER_10_193 ();
 fill_1 FILLER_10_195 ();
 decap_12 FILLER_10_197 ();
 decap_12 FILLER_10_209 ();
 decap_12 FILLER_10_221 ();
 decap_12 FILLER_10_233 ();
 fill_4 FILLER_10_245 ();
 fill_2 FILLER_10_249 ();
 fill_1 FILLER_10_251 ();
 decap_12 FILLER_10_253 ();
 decap_12 FILLER_10_265 ();
 decap_12 FILLER_10_277 ();
 decap_12 FILLER_10_289 ();
 fill_4 FILLER_10_301 ();
 fill_2 FILLER_10_305 ();
 fill_1 FILLER_10_307 ();
 decap_12 FILLER_10_309 ();
 decap_12 FILLER_10_321 ();
 decap_12 FILLER_10_333 ();
 decap_12 FILLER_10_345 ();
 fill_4 FILLER_10_357 ();
 fill_2 FILLER_10_361 ();
 fill_1 FILLER_10_363 ();
 decap_12 FILLER_10_365 ();
 decap_12 FILLER_10_377 ();
 decap_12 FILLER_10_389 ();
 decap_12 FILLER_10_401 ();
 fill_4 FILLER_10_413 ();
 fill_2 FILLER_10_417 ();
 fill_1 FILLER_10_419 ();
 decap_12 FILLER_10_421 ();
 decap_12 FILLER_10_433 ();
 decap_12 FILLER_10_445 ();
 decap_12 FILLER_10_457 ();
 fill_4 FILLER_10_469 ();
 fill_2 FILLER_10_473 ();
 fill_1 FILLER_10_475 ();
 decap_12 FILLER_10_477 ();
 decap_12 FILLER_10_489 ();
 decap_12 FILLER_10_501 ();
 decap_12 FILLER_10_513 ();
 fill_4 FILLER_10_525 ();
 fill_2 FILLER_10_529 ();
 fill_1 FILLER_10_531 ();
 decap_12 FILLER_10_533 ();
 decap_12 FILLER_10_545 ();
 decap_12 FILLER_10_557 ();
 decap_12 FILLER_10_569 ();
 fill_4 FILLER_10_581 ();
 fill_2 FILLER_10_585 ();
 fill_1 FILLER_10_587 ();
 decap_12 FILLER_10_589 ();
 decap_12 FILLER_10_601 ();
 decap_12 FILLER_10_613 ();
 decap_12 FILLER_11_3 ();
 decap_12 FILLER_11_15 ();
 decap_12 FILLER_11_27 ();
 decap_12 FILLER_11_39 ();
 fill_4 FILLER_11_51 ();
 fill_1 FILLER_11_55 ();
 decap_12 FILLER_11_57 ();
 decap_12 FILLER_11_69 ();
 decap_12 FILLER_11_81 ();
 decap_12 FILLER_11_93 ();
 fill_4 FILLER_11_105 ();
 fill_2 FILLER_11_109 ();
 fill_1 FILLER_11_111 ();
 decap_12 FILLER_11_113 ();
 decap_12 FILLER_11_125 ();
 decap_12 FILLER_11_137 ();
 decap_12 FILLER_11_149 ();
 fill_4 FILLER_11_161 ();
 fill_2 FILLER_11_165 ();
 fill_1 FILLER_11_167 ();
 decap_12 FILLER_11_169 ();
 decap_12 FILLER_11_181 ();
 decap_12 FILLER_11_193 ();
 decap_12 FILLER_11_205 ();
 fill_4 FILLER_11_217 ();
 fill_2 FILLER_11_221 ();
 fill_1 FILLER_11_223 ();
 decap_12 FILLER_11_225 ();
 decap_12 FILLER_11_237 ();
 decap_12 FILLER_11_249 ();
 decap_12 FILLER_11_261 ();
 fill_4 FILLER_11_273 ();
 fill_2 FILLER_11_277 ();
 fill_1 FILLER_11_279 ();
 decap_12 FILLER_11_281 ();
 decap_12 FILLER_11_293 ();
 decap_12 FILLER_11_305 ();
 decap_12 FILLER_11_317 ();
 fill_4 FILLER_11_329 ();
 fill_2 FILLER_11_333 ();
 fill_1 FILLER_11_335 ();
 decap_12 FILLER_11_337 ();
 decap_12 FILLER_11_349 ();
 decap_12 FILLER_11_361 ();
 decap_12 FILLER_11_373 ();
 fill_4 FILLER_11_385 ();
 fill_2 FILLER_11_389 ();
 fill_1 FILLER_11_391 ();
 decap_12 FILLER_11_393 ();
 decap_12 FILLER_11_405 ();
 decap_12 FILLER_11_417 ();
 decap_12 FILLER_11_429 ();
 fill_4 FILLER_11_441 ();
 fill_2 FILLER_11_445 ();
 fill_1 FILLER_11_447 ();
 decap_12 FILLER_11_449 ();
 decap_12 FILLER_11_461 ();
 decap_12 FILLER_11_473 ();
 decap_12 FILLER_11_485 ();
 fill_4 FILLER_11_497 ();
 fill_2 FILLER_11_501 ();
 fill_1 FILLER_11_503 ();
 decap_12 FILLER_11_505 ();
 decap_12 FILLER_11_517 ();
 decap_12 FILLER_11_529 ();
 decap_12 FILLER_11_541 ();
 fill_4 FILLER_11_553 ();
 fill_2 FILLER_11_557 ();
 fill_1 FILLER_11_559 ();
 decap_12 FILLER_11_561 ();
 decap_12 FILLER_11_573 ();
 decap_12 FILLER_11_585 ();
 decap_12 FILLER_11_597 ();
 fill_4 FILLER_11_609 ();
 fill_2 FILLER_11_613 ();
 fill_1 FILLER_11_615 ();
 fill_8 FILLER_11_617 ();
 decap_12 FILLER_12_3 ();
 decap_12 FILLER_12_15 ();
 fill_1 FILLER_12_27 ();
 decap_12 FILLER_12_29 ();
 decap_12 FILLER_12_41 ();
 decap_12 FILLER_12_53 ();
 decap_12 FILLER_12_65 ();
 fill_4 FILLER_12_77 ();
 fill_2 FILLER_12_81 ();
 fill_1 FILLER_12_83 ();
 decap_12 FILLER_12_85 ();
 decap_12 FILLER_12_97 ();
 decap_12 FILLER_12_109 ();
 decap_12 FILLER_12_121 ();
 fill_4 FILLER_12_133 ();
 fill_2 FILLER_12_137 ();
 fill_1 FILLER_12_139 ();
 decap_12 FILLER_12_141 ();
 decap_12 FILLER_12_153 ();
 decap_12 FILLER_12_165 ();
 decap_12 FILLER_12_177 ();
 fill_4 FILLER_12_189 ();
 fill_2 FILLER_12_193 ();
 fill_1 FILLER_12_195 ();
 decap_12 FILLER_12_197 ();
 decap_12 FILLER_12_209 ();
 decap_12 FILLER_12_221 ();
 decap_12 FILLER_12_233 ();
 fill_4 FILLER_12_245 ();
 fill_2 FILLER_12_249 ();
 fill_1 FILLER_12_251 ();
 decap_12 FILLER_12_253 ();
 decap_12 FILLER_12_265 ();
 decap_12 FILLER_12_277 ();
 decap_12 FILLER_12_289 ();
 fill_4 FILLER_12_301 ();
 fill_2 FILLER_12_305 ();
 fill_1 FILLER_12_307 ();
 decap_12 FILLER_12_309 ();
 decap_12 FILLER_12_321 ();
 decap_12 FILLER_12_333 ();
 decap_12 FILLER_12_345 ();
 fill_4 FILLER_12_357 ();
 fill_2 FILLER_12_361 ();
 fill_1 FILLER_12_363 ();
 decap_12 FILLER_12_365 ();
 decap_12 FILLER_12_377 ();
 decap_12 FILLER_12_389 ();
 decap_12 FILLER_12_401 ();
 fill_4 FILLER_12_413 ();
 fill_2 FILLER_12_417 ();
 fill_1 FILLER_12_419 ();
 decap_12 FILLER_12_421 ();
 decap_12 FILLER_12_433 ();
 decap_12 FILLER_12_445 ();
 decap_12 FILLER_12_457 ();
 fill_4 FILLER_12_469 ();
 fill_2 FILLER_12_473 ();
 fill_1 FILLER_12_475 ();
 decap_12 FILLER_12_477 ();
 decap_12 FILLER_12_489 ();
 decap_12 FILLER_12_501 ();
 decap_12 FILLER_12_513 ();
 fill_4 FILLER_12_525 ();
 fill_2 FILLER_12_529 ();
 fill_1 FILLER_12_531 ();
 decap_12 FILLER_12_533 ();
 decap_12 FILLER_12_545 ();
 decap_12 FILLER_12_557 ();
 decap_12 FILLER_12_569 ();
 fill_4 FILLER_12_581 ();
 fill_2 FILLER_12_585 ();
 fill_1 FILLER_12_587 ();
 decap_12 FILLER_12_589 ();
 decap_12 FILLER_12_601 ();
 decap_12 FILLER_12_613 ();
 decap_12 FILLER_13_3 ();
 decap_12 FILLER_13_15 ();
 decap_12 FILLER_13_27 ();
 decap_12 FILLER_13_39 ();
 fill_4 FILLER_13_51 ();
 fill_1 FILLER_13_55 ();
 decap_12 FILLER_13_57 ();
 decap_12 FILLER_13_69 ();
 decap_12 FILLER_13_81 ();
 decap_12 FILLER_13_93 ();
 fill_4 FILLER_13_105 ();
 fill_2 FILLER_13_109 ();
 fill_1 FILLER_13_111 ();
 decap_12 FILLER_13_113 ();
 decap_12 FILLER_13_125 ();
 decap_12 FILLER_13_137 ();
 decap_12 FILLER_13_149 ();
 fill_4 FILLER_13_161 ();
 fill_2 FILLER_13_165 ();
 fill_1 FILLER_13_167 ();
 decap_12 FILLER_13_169 ();
 decap_12 FILLER_13_181 ();
 decap_12 FILLER_13_193 ();
 decap_12 FILLER_13_205 ();
 fill_4 FILLER_13_217 ();
 fill_2 FILLER_13_221 ();
 fill_1 FILLER_13_223 ();
 decap_12 FILLER_13_225 ();
 decap_12 FILLER_13_237 ();
 decap_12 FILLER_13_249 ();
 decap_12 FILLER_13_261 ();
 fill_4 FILLER_13_273 ();
 fill_2 FILLER_13_277 ();
 fill_1 FILLER_13_279 ();
 decap_12 FILLER_13_281 ();
 decap_12 FILLER_13_293 ();
 decap_12 FILLER_13_305 ();
 decap_12 FILLER_13_317 ();
 fill_4 FILLER_13_329 ();
 fill_2 FILLER_13_333 ();
 fill_1 FILLER_13_335 ();
 decap_12 FILLER_13_337 ();
 decap_12 FILLER_13_349 ();
 decap_12 FILLER_13_361 ();
 decap_12 FILLER_13_373 ();
 fill_4 FILLER_13_385 ();
 fill_2 FILLER_13_389 ();
 fill_1 FILLER_13_391 ();
 decap_12 FILLER_13_393 ();
 decap_12 FILLER_13_405 ();
 decap_12 FILLER_13_417 ();
 decap_12 FILLER_13_429 ();
 fill_4 FILLER_13_441 ();
 fill_2 FILLER_13_445 ();
 fill_1 FILLER_13_447 ();
 decap_12 FILLER_13_449 ();
 decap_12 FILLER_13_461 ();
 decap_12 FILLER_13_473 ();
 decap_12 FILLER_13_485 ();
 fill_4 FILLER_13_497 ();
 fill_2 FILLER_13_501 ();
 fill_1 FILLER_13_503 ();
 decap_12 FILLER_13_505 ();
 decap_12 FILLER_13_517 ();
 decap_12 FILLER_13_529 ();
 decap_12 FILLER_13_541 ();
 fill_4 FILLER_13_553 ();
 fill_2 FILLER_13_557 ();
 fill_1 FILLER_13_559 ();
 decap_12 FILLER_13_561 ();
 decap_12 FILLER_13_573 ();
 decap_12 FILLER_13_585 ();
 decap_12 FILLER_13_597 ();
 fill_4 FILLER_13_609 ();
 fill_2 FILLER_13_613 ();
 fill_1 FILLER_13_615 ();
 fill_8 FILLER_13_617 ();
 decap_12 FILLER_14_3 ();
 decap_12 FILLER_14_15 ();
 fill_1 FILLER_14_27 ();
 decap_12 FILLER_14_29 ();
 decap_12 FILLER_14_41 ();
 decap_12 FILLER_14_53 ();
 decap_12 FILLER_14_65 ();
 fill_4 FILLER_14_77 ();
 fill_2 FILLER_14_81 ();
 fill_1 FILLER_14_83 ();
 decap_12 FILLER_14_85 ();
 decap_12 FILLER_14_97 ();
 decap_12 FILLER_14_109 ();
 decap_12 FILLER_14_121 ();
 fill_4 FILLER_14_133 ();
 fill_2 FILLER_14_137 ();
 fill_1 FILLER_14_139 ();
 decap_12 FILLER_14_141 ();
 decap_12 FILLER_14_153 ();
 decap_12 FILLER_14_165 ();
 decap_12 FILLER_14_177 ();
 fill_4 FILLER_14_189 ();
 fill_2 FILLER_14_193 ();
 fill_1 FILLER_14_195 ();
 decap_12 FILLER_14_197 ();
 decap_12 FILLER_14_209 ();
 decap_12 FILLER_14_221 ();
 decap_12 FILLER_14_233 ();
 fill_4 FILLER_14_245 ();
 fill_2 FILLER_14_249 ();
 fill_1 FILLER_14_251 ();
 decap_12 FILLER_14_253 ();
 decap_12 FILLER_14_265 ();
 decap_12 FILLER_14_277 ();
 decap_12 FILLER_14_289 ();
 fill_4 FILLER_14_301 ();
 fill_2 FILLER_14_305 ();
 fill_1 FILLER_14_307 ();
 decap_12 FILLER_14_309 ();
 decap_12 FILLER_14_321 ();
 decap_12 FILLER_14_333 ();
 decap_12 FILLER_14_345 ();
 fill_4 FILLER_14_357 ();
 fill_2 FILLER_14_361 ();
 fill_1 FILLER_14_363 ();
 decap_12 FILLER_14_365 ();
 decap_12 FILLER_14_377 ();
 decap_12 FILLER_14_389 ();
 decap_12 FILLER_14_401 ();
 fill_4 FILLER_14_413 ();
 fill_2 FILLER_14_417 ();
 fill_1 FILLER_14_419 ();
 decap_12 FILLER_14_421 ();
 decap_12 FILLER_14_433 ();
 decap_12 FILLER_14_445 ();
 decap_12 FILLER_14_457 ();
 fill_4 FILLER_14_469 ();
 fill_2 FILLER_14_473 ();
 fill_1 FILLER_14_475 ();
 decap_12 FILLER_14_477 ();
 decap_12 FILLER_14_489 ();
 decap_12 FILLER_14_501 ();
 decap_12 FILLER_14_513 ();
 fill_4 FILLER_14_525 ();
 fill_2 FILLER_14_529 ();
 fill_1 FILLER_14_531 ();
 decap_12 FILLER_14_533 ();
 decap_12 FILLER_14_545 ();
 decap_12 FILLER_14_557 ();
 decap_12 FILLER_14_569 ();
 fill_4 FILLER_14_581 ();
 fill_2 FILLER_14_585 ();
 fill_1 FILLER_14_587 ();
 decap_12 FILLER_14_589 ();
 decap_12 FILLER_14_601 ();
 decap_12 FILLER_14_613 ();
 decap_12 FILLER_15_3 ();
 decap_12 FILLER_15_15 ();
 decap_12 FILLER_15_27 ();
 decap_12 FILLER_15_39 ();
 fill_4 FILLER_15_51 ();
 fill_1 FILLER_15_55 ();
 decap_12 FILLER_15_57 ();
 decap_12 FILLER_15_69 ();
 decap_12 FILLER_15_81 ();
 decap_12 FILLER_15_93 ();
 fill_4 FILLER_15_105 ();
 fill_2 FILLER_15_109 ();
 fill_1 FILLER_15_111 ();
 decap_12 FILLER_15_113 ();
 decap_12 FILLER_15_125 ();
 decap_12 FILLER_15_137 ();
 decap_12 FILLER_15_149 ();
 fill_4 FILLER_15_161 ();
 fill_2 FILLER_15_165 ();
 fill_1 FILLER_15_167 ();
 decap_12 FILLER_15_169 ();
 decap_12 FILLER_15_181 ();
 decap_12 FILLER_15_193 ();
 decap_12 FILLER_15_205 ();
 fill_4 FILLER_15_217 ();
 fill_2 FILLER_15_221 ();
 fill_1 FILLER_15_223 ();
 decap_12 FILLER_15_225 ();
 decap_12 FILLER_15_237 ();
 decap_12 FILLER_15_249 ();
 decap_12 FILLER_15_261 ();
 fill_4 FILLER_15_273 ();
 fill_2 FILLER_15_277 ();
 fill_1 FILLER_15_279 ();
 decap_12 FILLER_15_281 ();
 decap_12 FILLER_15_293 ();
 decap_12 FILLER_15_305 ();
 decap_12 FILLER_15_317 ();
 fill_4 FILLER_15_329 ();
 fill_2 FILLER_15_333 ();
 fill_1 FILLER_15_335 ();
 decap_12 FILLER_15_337 ();
 decap_12 FILLER_15_349 ();
 decap_12 FILLER_15_361 ();
 decap_12 FILLER_15_373 ();
 fill_4 FILLER_15_385 ();
 fill_2 FILLER_15_389 ();
 fill_1 FILLER_15_391 ();
 decap_12 FILLER_15_393 ();
 decap_12 FILLER_15_405 ();
 decap_12 FILLER_15_417 ();
 decap_12 FILLER_15_429 ();
 fill_4 FILLER_15_441 ();
 fill_2 FILLER_15_445 ();
 fill_1 FILLER_15_447 ();
 decap_12 FILLER_15_449 ();
 decap_12 FILLER_15_461 ();
 decap_12 FILLER_15_473 ();
 decap_12 FILLER_15_485 ();
 fill_4 FILLER_15_497 ();
 fill_2 FILLER_15_501 ();
 fill_1 FILLER_15_503 ();
 decap_12 FILLER_15_505 ();
 decap_12 FILLER_15_517 ();
 decap_12 FILLER_15_529 ();
 decap_12 FILLER_15_541 ();
 fill_4 FILLER_15_553 ();
 fill_2 FILLER_15_557 ();
 fill_1 FILLER_15_559 ();
 decap_12 FILLER_15_561 ();
 decap_12 FILLER_15_573 ();
 decap_12 FILLER_15_585 ();
 decap_12 FILLER_15_597 ();
 fill_4 FILLER_15_609 ();
 fill_2 FILLER_15_613 ();
 fill_1 FILLER_15_615 ();
 fill_8 FILLER_15_617 ();
 decap_12 FILLER_16_3 ();
 decap_12 FILLER_16_15 ();
 fill_1 FILLER_16_27 ();
 decap_12 FILLER_16_29 ();
 decap_12 FILLER_16_41 ();
 decap_12 FILLER_16_53 ();
 decap_12 FILLER_16_65 ();
 fill_4 FILLER_16_77 ();
 fill_2 FILLER_16_81 ();
 fill_1 FILLER_16_83 ();
 decap_12 FILLER_16_85 ();
 decap_12 FILLER_16_97 ();
 decap_12 FILLER_16_109 ();
 decap_12 FILLER_16_121 ();
 fill_4 FILLER_16_133 ();
 fill_2 FILLER_16_137 ();
 fill_1 FILLER_16_139 ();
 decap_12 FILLER_16_141 ();
 decap_12 FILLER_16_153 ();
 decap_12 FILLER_16_165 ();
 decap_12 FILLER_16_177 ();
 fill_4 FILLER_16_189 ();
 fill_2 FILLER_16_193 ();
 fill_1 FILLER_16_195 ();
 decap_12 FILLER_16_197 ();
 decap_12 FILLER_16_209 ();
 decap_12 FILLER_16_221 ();
 decap_12 FILLER_16_233 ();
 fill_4 FILLER_16_245 ();
 fill_2 FILLER_16_249 ();
 fill_1 FILLER_16_251 ();
 decap_12 FILLER_16_253 ();
 decap_12 FILLER_16_265 ();
 decap_12 FILLER_16_277 ();
 decap_12 FILLER_16_289 ();
 fill_4 FILLER_16_301 ();
 fill_2 FILLER_16_305 ();
 fill_1 FILLER_16_307 ();
 decap_12 FILLER_16_309 ();
 decap_12 FILLER_16_321 ();
 decap_12 FILLER_16_333 ();
 decap_12 FILLER_16_345 ();
 fill_4 FILLER_16_357 ();
 fill_2 FILLER_16_361 ();
 fill_1 FILLER_16_363 ();
 decap_12 FILLER_16_365 ();
 decap_12 FILLER_16_377 ();
 decap_12 FILLER_16_389 ();
 decap_12 FILLER_16_401 ();
 fill_4 FILLER_16_413 ();
 fill_2 FILLER_16_417 ();
 fill_1 FILLER_16_419 ();
 decap_12 FILLER_16_421 ();
 decap_12 FILLER_16_433 ();
 decap_12 FILLER_16_445 ();
 decap_12 FILLER_16_457 ();
 fill_4 FILLER_16_469 ();
 fill_2 FILLER_16_473 ();
 fill_1 FILLER_16_475 ();
 decap_12 FILLER_16_477 ();
 decap_12 FILLER_16_489 ();
 decap_12 FILLER_16_501 ();
 decap_12 FILLER_16_513 ();
 fill_4 FILLER_16_525 ();
 fill_2 FILLER_16_529 ();
 fill_1 FILLER_16_531 ();
 decap_12 FILLER_16_533 ();
 decap_12 FILLER_16_545 ();
 decap_12 FILLER_16_557 ();
 decap_12 FILLER_16_569 ();
 fill_4 FILLER_16_581 ();
 fill_2 FILLER_16_585 ();
 fill_1 FILLER_16_587 ();
 decap_12 FILLER_16_589 ();
 decap_12 FILLER_16_601 ();
 decap_12 FILLER_16_613 ();
 decap_12 FILLER_17_3 ();
 decap_12 FILLER_17_15 ();
 decap_12 FILLER_17_27 ();
 decap_12 FILLER_17_39 ();
 fill_4 FILLER_17_51 ();
 fill_1 FILLER_17_55 ();
 decap_12 FILLER_17_57 ();
 decap_12 FILLER_17_69 ();
 decap_12 FILLER_17_81 ();
 decap_12 FILLER_17_93 ();
 fill_4 FILLER_17_105 ();
 fill_2 FILLER_17_109 ();
 fill_1 FILLER_17_111 ();
 decap_12 FILLER_17_113 ();
 decap_12 FILLER_17_125 ();
 decap_12 FILLER_17_137 ();
 decap_12 FILLER_17_149 ();
 fill_4 FILLER_17_161 ();
 fill_2 FILLER_17_165 ();
 fill_1 FILLER_17_167 ();
 decap_12 FILLER_17_169 ();
 decap_12 FILLER_17_181 ();
 decap_12 FILLER_17_193 ();
 decap_12 FILLER_17_205 ();
 fill_4 FILLER_17_217 ();
 fill_2 FILLER_17_221 ();
 fill_1 FILLER_17_223 ();
 decap_12 FILLER_17_225 ();
 decap_12 FILLER_17_237 ();
 decap_12 FILLER_17_249 ();
 decap_12 FILLER_17_261 ();
 fill_4 FILLER_17_273 ();
 fill_2 FILLER_17_277 ();
 fill_1 FILLER_17_279 ();
 decap_12 FILLER_17_281 ();
 decap_12 FILLER_17_293 ();
 decap_12 FILLER_17_305 ();
 decap_12 FILLER_17_317 ();
 fill_4 FILLER_17_329 ();
 fill_2 FILLER_17_333 ();
 fill_1 FILLER_17_335 ();
 decap_12 FILLER_17_337 ();
 decap_12 FILLER_17_349 ();
 decap_12 FILLER_17_361 ();
 decap_12 FILLER_17_373 ();
 fill_4 FILLER_17_385 ();
 fill_2 FILLER_17_389 ();
 fill_1 FILLER_17_391 ();
 decap_12 FILLER_17_393 ();
 decap_12 FILLER_17_405 ();
 decap_12 FILLER_17_417 ();
 decap_12 FILLER_17_429 ();
 fill_4 FILLER_17_441 ();
 fill_2 FILLER_17_445 ();
 fill_1 FILLER_17_447 ();
 decap_12 FILLER_17_449 ();
 decap_12 FILLER_17_461 ();
 decap_12 FILLER_17_473 ();
 decap_12 FILLER_17_485 ();
 fill_4 FILLER_17_497 ();
 fill_2 FILLER_17_501 ();
 fill_1 FILLER_17_503 ();
 decap_12 FILLER_17_505 ();
 decap_12 FILLER_17_517 ();
 decap_12 FILLER_17_529 ();
 decap_12 FILLER_17_541 ();
 fill_4 FILLER_17_553 ();
 fill_2 FILLER_17_557 ();
 fill_1 FILLER_17_559 ();
 decap_12 FILLER_17_561 ();
 decap_12 FILLER_17_573 ();
 decap_12 FILLER_17_585 ();
 decap_12 FILLER_17_597 ();
 fill_4 FILLER_17_609 ();
 fill_2 FILLER_17_613 ();
 fill_1 FILLER_17_615 ();
 fill_8 FILLER_17_617 ();
 decap_12 FILLER_18_3 ();
 decap_12 FILLER_18_15 ();
 fill_1 FILLER_18_27 ();
 decap_12 FILLER_18_29 ();
 decap_12 FILLER_18_41 ();
 decap_12 FILLER_18_53 ();
 decap_12 FILLER_18_65 ();
 fill_4 FILLER_18_77 ();
 fill_2 FILLER_18_81 ();
 fill_1 FILLER_18_83 ();
 decap_12 FILLER_18_85 ();
 decap_12 FILLER_18_97 ();
 decap_12 FILLER_18_109 ();
 decap_12 FILLER_18_121 ();
 fill_4 FILLER_18_133 ();
 fill_2 FILLER_18_137 ();
 fill_1 FILLER_18_139 ();
 decap_12 FILLER_18_141 ();
 decap_12 FILLER_18_153 ();
 decap_12 FILLER_18_165 ();
 decap_12 FILLER_18_177 ();
 fill_4 FILLER_18_189 ();
 fill_2 FILLER_18_193 ();
 fill_1 FILLER_18_195 ();
 decap_12 FILLER_18_197 ();
 decap_12 FILLER_18_209 ();
 decap_12 FILLER_18_221 ();
 decap_12 FILLER_18_233 ();
 fill_4 FILLER_18_245 ();
 fill_2 FILLER_18_249 ();
 fill_1 FILLER_18_251 ();
 decap_12 FILLER_18_253 ();
 decap_12 FILLER_18_265 ();
 decap_12 FILLER_18_277 ();
 decap_12 FILLER_18_289 ();
 fill_4 FILLER_18_301 ();
 fill_2 FILLER_18_305 ();
 fill_1 FILLER_18_307 ();
 decap_12 FILLER_18_309 ();
 decap_12 FILLER_18_321 ();
 decap_12 FILLER_18_333 ();
 decap_12 FILLER_18_345 ();
 fill_4 FILLER_18_357 ();
 fill_2 FILLER_18_361 ();
 fill_1 FILLER_18_363 ();
 decap_12 FILLER_18_365 ();
 decap_12 FILLER_18_377 ();
 decap_12 FILLER_18_389 ();
 decap_12 FILLER_18_401 ();
 fill_4 FILLER_18_413 ();
 fill_2 FILLER_18_417 ();
 fill_1 FILLER_18_419 ();
 decap_12 FILLER_18_421 ();
 decap_12 FILLER_18_433 ();
 decap_12 FILLER_18_445 ();
 decap_12 FILLER_18_457 ();
 fill_4 FILLER_18_469 ();
 fill_2 FILLER_18_473 ();
 fill_1 FILLER_18_475 ();
 decap_12 FILLER_18_477 ();
 decap_12 FILLER_18_489 ();
 decap_12 FILLER_18_501 ();
 decap_12 FILLER_18_513 ();
 fill_4 FILLER_18_525 ();
 fill_2 FILLER_18_529 ();
 fill_1 FILLER_18_531 ();
 decap_12 FILLER_18_533 ();
 decap_12 FILLER_18_545 ();
 decap_12 FILLER_18_557 ();
 decap_12 FILLER_18_569 ();
 fill_4 FILLER_18_581 ();
 fill_2 FILLER_18_585 ();
 fill_1 FILLER_18_587 ();
 decap_12 FILLER_18_589 ();
 decap_12 FILLER_18_601 ();
 decap_12 FILLER_18_613 ();
 decap_12 FILLER_19_3 ();
 decap_12 FILLER_19_15 ();
 decap_12 FILLER_19_27 ();
 decap_12 FILLER_19_39 ();
 fill_4 FILLER_19_51 ();
 fill_1 FILLER_19_55 ();
 decap_12 FILLER_19_57 ();
 decap_12 FILLER_19_69 ();
 decap_12 FILLER_19_81 ();
 decap_12 FILLER_19_93 ();
 fill_4 FILLER_19_105 ();
 fill_2 FILLER_19_109 ();
 fill_1 FILLER_19_111 ();
 decap_12 FILLER_19_113 ();
 decap_12 FILLER_19_125 ();
 decap_12 FILLER_19_137 ();
 decap_12 FILLER_19_149 ();
 fill_4 FILLER_19_161 ();
 fill_2 FILLER_19_165 ();
 fill_1 FILLER_19_167 ();
 decap_12 FILLER_19_169 ();
 decap_12 FILLER_19_181 ();
 decap_12 FILLER_19_193 ();
 decap_12 FILLER_19_205 ();
 fill_4 FILLER_19_217 ();
 fill_2 FILLER_19_221 ();
 fill_1 FILLER_19_223 ();
 decap_12 FILLER_19_225 ();
 decap_12 FILLER_19_237 ();
 decap_12 FILLER_19_249 ();
 decap_12 FILLER_19_261 ();
 fill_4 FILLER_19_273 ();
 fill_2 FILLER_19_277 ();
 fill_1 FILLER_19_279 ();
 decap_12 FILLER_19_281 ();
 decap_12 FILLER_19_293 ();
 decap_12 FILLER_19_305 ();
 decap_12 FILLER_19_317 ();
 fill_4 FILLER_19_329 ();
 fill_2 FILLER_19_333 ();
 fill_1 FILLER_19_335 ();
 decap_12 FILLER_19_337 ();
 decap_12 FILLER_19_349 ();
 decap_12 FILLER_19_361 ();
 decap_12 FILLER_19_373 ();
 fill_4 FILLER_19_385 ();
 fill_2 FILLER_19_389 ();
 fill_1 FILLER_19_391 ();
 decap_12 FILLER_19_393 ();
 decap_12 FILLER_19_405 ();
 decap_12 FILLER_19_417 ();
 decap_12 FILLER_19_429 ();
 fill_4 FILLER_19_441 ();
 fill_2 FILLER_19_445 ();
 fill_1 FILLER_19_447 ();
 decap_12 FILLER_19_449 ();
 decap_12 FILLER_19_461 ();
 decap_12 FILLER_19_473 ();
 decap_12 FILLER_19_485 ();
 fill_4 FILLER_19_497 ();
 fill_2 FILLER_19_501 ();
 fill_1 FILLER_19_503 ();
 decap_12 FILLER_19_505 ();
 decap_12 FILLER_19_517 ();
 decap_12 FILLER_19_529 ();
 decap_12 FILLER_19_541 ();
 fill_4 FILLER_19_553 ();
 fill_2 FILLER_19_557 ();
 fill_1 FILLER_19_559 ();
 decap_12 FILLER_19_561 ();
 decap_12 FILLER_19_573 ();
 decap_12 FILLER_19_585 ();
 decap_12 FILLER_19_597 ();
 fill_4 FILLER_19_609 ();
 fill_2 FILLER_19_613 ();
 fill_1 FILLER_19_615 ();
 fill_8 FILLER_19_617 ();
 decap_12 FILLER_20_3 ();
 decap_12 FILLER_20_15 ();
 fill_1 FILLER_20_27 ();
 decap_12 FILLER_20_29 ();
 decap_12 FILLER_20_41 ();
 decap_12 FILLER_20_53 ();
 decap_12 FILLER_20_65 ();
 fill_4 FILLER_20_77 ();
 fill_2 FILLER_20_81 ();
 fill_1 FILLER_20_83 ();
 decap_12 FILLER_20_85 ();
 decap_12 FILLER_20_97 ();
 decap_12 FILLER_20_109 ();
 decap_12 FILLER_20_121 ();
 fill_4 FILLER_20_133 ();
 fill_2 FILLER_20_137 ();
 fill_1 FILLER_20_139 ();
 decap_12 FILLER_20_141 ();
 decap_12 FILLER_20_153 ();
 decap_12 FILLER_20_165 ();
 decap_12 FILLER_20_177 ();
 fill_4 FILLER_20_189 ();
 fill_2 FILLER_20_193 ();
 fill_1 FILLER_20_195 ();
 decap_12 FILLER_20_197 ();
 decap_12 FILLER_20_209 ();
 decap_12 FILLER_20_221 ();
 decap_12 FILLER_20_233 ();
 fill_4 FILLER_20_245 ();
 fill_2 FILLER_20_249 ();
 fill_1 FILLER_20_251 ();
 decap_12 FILLER_20_253 ();
 decap_12 FILLER_20_265 ();
 decap_12 FILLER_20_277 ();
 decap_12 FILLER_20_289 ();
 fill_4 FILLER_20_301 ();
 fill_2 FILLER_20_305 ();
 fill_1 FILLER_20_307 ();
 decap_12 FILLER_20_309 ();
 decap_12 FILLER_20_321 ();
 decap_12 FILLER_20_333 ();
 decap_12 FILLER_20_345 ();
 fill_4 FILLER_20_357 ();
 fill_2 FILLER_20_361 ();
 fill_1 FILLER_20_363 ();
 decap_12 FILLER_20_365 ();
 decap_12 FILLER_20_377 ();
 decap_12 FILLER_20_389 ();
 decap_12 FILLER_20_401 ();
 fill_4 FILLER_20_413 ();
 fill_2 FILLER_20_417 ();
 fill_1 FILLER_20_419 ();
 decap_12 FILLER_20_421 ();
 decap_12 FILLER_20_433 ();
 decap_12 FILLER_20_445 ();
 decap_12 FILLER_20_457 ();
 fill_4 FILLER_20_469 ();
 fill_2 FILLER_20_473 ();
 fill_1 FILLER_20_475 ();
 decap_12 FILLER_20_477 ();
 decap_12 FILLER_20_489 ();
 decap_12 FILLER_20_501 ();
 decap_12 FILLER_20_513 ();
 fill_4 FILLER_20_525 ();
 fill_2 FILLER_20_529 ();
 fill_1 FILLER_20_531 ();
 decap_12 FILLER_20_533 ();
 decap_12 FILLER_20_545 ();
 decap_12 FILLER_20_557 ();
 decap_12 FILLER_20_569 ();
 fill_4 FILLER_20_581 ();
 fill_2 FILLER_20_585 ();
 fill_1 FILLER_20_587 ();
 decap_12 FILLER_20_589 ();
 decap_12 FILLER_20_601 ();
 decap_12 FILLER_20_613 ();
 decap_12 FILLER_21_3 ();
 decap_12 FILLER_21_15 ();
 decap_12 FILLER_21_27 ();
 decap_12 FILLER_21_39 ();
 fill_4 FILLER_21_51 ();
 fill_1 FILLER_21_55 ();
 decap_12 FILLER_21_57 ();
 decap_12 FILLER_21_69 ();
 decap_12 FILLER_21_81 ();
 decap_12 FILLER_21_93 ();
 fill_4 FILLER_21_105 ();
 fill_2 FILLER_21_109 ();
 fill_1 FILLER_21_111 ();
 decap_12 FILLER_21_113 ();
 decap_12 FILLER_21_125 ();
 decap_12 FILLER_21_137 ();
 decap_12 FILLER_21_149 ();
 fill_4 FILLER_21_161 ();
 fill_2 FILLER_21_165 ();
 fill_1 FILLER_21_167 ();
 decap_12 FILLER_21_169 ();
 decap_12 FILLER_21_181 ();
 decap_12 FILLER_21_193 ();
 decap_12 FILLER_21_205 ();
 fill_4 FILLER_21_217 ();
 fill_2 FILLER_21_221 ();
 fill_1 FILLER_21_223 ();
 decap_12 FILLER_21_225 ();
 decap_12 FILLER_21_237 ();
 decap_12 FILLER_21_249 ();
 decap_12 FILLER_21_261 ();
 fill_4 FILLER_21_273 ();
 fill_2 FILLER_21_277 ();
 fill_1 FILLER_21_279 ();
 decap_12 FILLER_21_281 ();
 decap_12 FILLER_21_293 ();
 decap_12 FILLER_21_305 ();
 decap_12 FILLER_21_317 ();
 fill_4 FILLER_21_329 ();
 fill_2 FILLER_21_333 ();
 fill_1 FILLER_21_335 ();
 decap_12 FILLER_21_337 ();
 decap_12 FILLER_21_349 ();
 decap_12 FILLER_21_361 ();
 decap_12 FILLER_21_373 ();
 fill_4 FILLER_21_385 ();
 fill_2 FILLER_21_389 ();
 fill_1 FILLER_21_391 ();
 decap_12 FILLER_21_393 ();
 decap_12 FILLER_21_405 ();
 decap_12 FILLER_21_417 ();
 decap_12 FILLER_21_429 ();
 fill_4 FILLER_21_441 ();
 fill_2 FILLER_21_445 ();
 fill_1 FILLER_21_447 ();
 decap_12 FILLER_21_449 ();
 decap_12 FILLER_21_461 ();
 decap_12 FILLER_21_473 ();
 decap_12 FILLER_21_485 ();
 fill_4 FILLER_21_497 ();
 fill_2 FILLER_21_501 ();
 fill_1 FILLER_21_503 ();
 decap_12 FILLER_21_505 ();
 decap_12 FILLER_21_517 ();
 decap_12 FILLER_21_529 ();
 decap_12 FILLER_21_541 ();
 fill_4 FILLER_21_553 ();
 fill_2 FILLER_21_557 ();
 fill_1 FILLER_21_559 ();
 decap_12 FILLER_21_561 ();
 decap_12 FILLER_21_573 ();
 decap_12 FILLER_21_585 ();
 decap_12 FILLER_21_597 ();
 fill_4 FILLER_21_609 ();
 fill_2 FILLER_21_613 ();
 fill_1 FILLER_21_615 ();
 fill_8 FILLER_21_617 ();
 decap_12 FILLER_22_3 ();
 decap_12 FILLER_22_15 ();
 fill_1 FILLER_22_27 ();
 decap_12 FILLER_22_29 ();
 decap_12 FILLER_22_41 ();
 decap_12 FILLER_22_53 ();
 decap_12 FILLER_22_65 ();
 fill_4 FILLER_22_77 ();
 fill_2 FILLER_22_81 ();
 fill_1 FILLER_22_83 ();
 decap_12 FILLER_22_85 ();
 decap_12 FILLER_22_97 ();
 decap_12 FILLER_22_109 ();
 decap_12 FILLER_22_121 ();
 fill_4 FILLER_22_133 ();
 fill_2 FILLER_22_137 ();
 fill_1 FILLER_22_139 ();
 decap_12 FILLER_22_141 ();
 decap_12 FILLER_22_153 ();
 decap_12 FILLER_22_165 ();
 decap_12 FILLER_22_177 ();
 fill_4 FILLER_22_189 ();
 fill_2 FILLER_22_193 ();
 fill_1 FILLER_22_195 ();
 decap_12 FILLER_22_197 ();
 decap_12 FILLER_22_209 ();
 decap_12 FILLER_22_221 ();
 decap_12 FILLER_22_233 ();
 fill_4 FILLER_22_245 ();
 fill_2 FILLER_22_249 ();
 fill_1 FILLER_22_251 ();
 decap_12 FILLER_22_253 ();
 decap_12 FILLER_22_265 ();
 decap_12 FILLER_22_277 ();
 decap_12 FILLER_22_289 ();
 fill_4 FILLER_22_301 ();
 fill_2 FILLER_22_305 ();
 fill_1 FILLER_22_307 ();
 decap_12 FILLER_22_309 ();
 decap_12 FILLER_22_321 ();
 decap_12 FILLER_22_333 ();
 decap_12 FILLER_22_345 ();
 fill_4 FILLER_22_357 ();
 fill_2 FILLER_22_361 ();
 fill_1 FILLER_22_363 ();
 decap_12 FILLER_22_365 ();
 decap_12 FILLER_22_377 ();
 decap_12 FILLER_22_389 ();
 decap_12 FILLER_22_401 ();
 fill_4 FILLER_22_413 ();
 fill_2 FILLER_22_417 ();
 fill_1 FILLER_22_419 ();
 decap_12 FILLER_22_421 ();
 decap_12 FILLER_22_433 ();
 decap_12 FILLER_22_445 ();
 decap_12 FILLER_22_457 ();
 fill_4 FILLER_22_469 ();
 fill_2 FILLER_22_473 ();
 fill_1 FILLER_22_475 ();
 decap_12 FILLER_22_477 ();
 decap_12 FILLER_22_489 ();
 decap_12 FILLER_22_501 ();
 decap_12 FILLER_22_513 ();
 fill_4 FILLER_22_525 ();
 fill_2 FILLER_22_529 ();
 fill_1 FILLER_22_531 ();
 decap_12 FILLER_22_533 ();
 decap_12 FILLER_22_545 ();
 decap_12 FILLER_22_557 ();
 decap_12 FILLER_22_569 ();
 fill_4 FILLER_22_581 ();
 fill_2 FILLER_22_585 ();
 fill_1 FILLER_22_587 ();
 decap_12 FILLER_22_589 ();
 decap_12 FILLER_22_601 ();
 decap_12 FILLER_22_613 ();
 decap_12 FILLER_23_3 ();
 decap_12 FILLER_23_15 ();
 decap_12 FILLER_23_27 ();
 decap_12 FILLER_23_39 ();
 fill_4 FILLER_23_51 ();
 fill_1 FILLER_23_55 ();
 decap_12 FILLER_23_57 ();
 decap_12 FILLER_23_69 ();
 decap_12 FILLER_23_81 ();
 decap_12 FILLER_23_93 ();
 fill_4 FILLER_23_105 ();
 fill_2 FILLER_23_109 ();
 fill_1 FILLER_23_111 ();
 decap_12 FILLER_23_113 ();
 decap_12 FILLER_23_125 ();
 decap_12 FILLER_23_137 ();
 decap_12 FILLER_23_149 ();
 fill_4 FILLER_23_161 ();
 fill_2 FILLER_23_165 ();
 fill_1 FILLER_23_167 ();
 decap_12 FILLER_23_169 ();
 decap_12 FILLER_23_181 ();
 decap_12 FILLER_23_193 ();
 decap_12 FILLER_23_205 ();
 fill_4 FILLER_23_217 ();
 fill_2 FILLER_23_221 ();
 fill_1 FILLER_23_223 ();
 decap_12 FILLER_23_225 ();
 decap_12 FILLER_23_237 ();
 decap_12 FILLER_23_249 ();
 decap_12 FILLER_23_261 ();
 fill_4 FILLER_23_273 ();
 fill_2 FILLER_23_277 ();
 fill_1 FILLER_23_279 ();
 decap_12 FILLER_23_281 ();
 decap_12 FILLER_23_293 ();
 decap_12 FILLER_23_305 ();
 decap_12 FILLER_23_317 ();
 fill_4 FILLER_23_329 ();
 fill_2 FILLER_23_333 ();
 fill_1 FILLER_23_335 ();
 decap_12 FILLER_23_337 ();
 decap_12 FILLER_23_349 ();
 decap_12 FILLER_23_361 ();
 decap_12 FILLER_23_373 ();
 fill_4 FILLER_23_385 ();
 fill_2 FILLER_23_389 ();
 fill_1 FILLER_23_391 ();
 decap_12 FILLER_23_393 ();
 decap_12 FILLER_23_405 ();
 decap_12 FILLER_23_417 ();
 decap_12 FILLER_23_429 ();
 fill_4 FILLER_23_441 ();
 fill_2 FILLER_23_445 ();
 fill_1 FILLER_23_447 ();
 decap_12 FILLER_23_449 ();
 decap_12 FILLER_23_461 ();
 decap_12 FILLER_23_473 ();
 decap_12 FILLER_23_485 ();
 fill_4 FILLER_23_497 ();
 fill_2 FILLER_23_501 ();
 fill_1 FILLER_23_503 ();
 decap_12 FILLER_23_505 ();
 decap_12 FILLER_23_517 ();
 decap_12 FILLER_23_529 ();
 decap_12 FILLER_23_541 ();
 fill_4 FILLER_23_553 ();
 fill_2 FILLER_23_557 ();
 fill_1 FILLER_23_559 ();
 decap_12 FILLER_23_561 ();
 decap_12 FILLER_23_573 ();
 decap_12 FILLER_23_585 ();
 decap_12 FILLER_23_597 ();
 fill_4 FILLER_23_609 ();
 fill_2 FILLER_23_613 ();
 fill_1 FILLER_23_615 ();
 fill_8 FILLER_23_617 ();
 decap_12 FILLER_24_3 ();
 decap_12 FILLER_24_15 ();
 fill_1 FILLER_24_27 ();
 decap_12 FILLER_24_29 ();
 decap_12 FILLER_24_41 ();
 decap_12 FILLER_24_53 ();
 decap_12 FILLER_24_65 ();
 fill_4 FILLER_24_77 ();
 fill_2 FILLER_24_81 ();
 fill_1 FILLER_24_83 ();
 decap_12 FILLER_24_85 ();
 decap_12 FILLER_24_97 ();
 decap_12 FILLER_24_109 ();
 decap_12 FILLER_24_121 ();
 fill_4 FILLER_24_133 ();
 fill_2 FILLER_24_137 ();
 fill_1 FILLER_24_139 ();
 decap_12 FILLER_24_141 ();
 decap_12 FILLER_24_153 ();
 decap_12 FILLER_24_165 ();
 decap_12 FILLER_24_177 ();
 fill_4 FILLER_24_189 ();
 fill_2 FILLER_24_193 ();
 fill_1 FILLER_24_195 ();
 decap_12 FILLER_24_197 ();
 decap_12 FILLER_24_209 ();
 decap_12 FILLER_24_221 ();
 decap_12 FILLER_24_233 ();
 fill_4 FILLER_24_245 ();
 fill_2 FILLER_24_249 ();
 fill_1 FILLER_24_251 ();
 decap_12 FILLER_24_253 ();
 decap_12 FILLER_24_265 ();
 decap_12 FILLER_24_277 ();
 decap_12 FILLER_24_289 ();
 fill_4 FILLER_24_301 ();
 fill_2 FILLER_24_305 ();
 fill_1 FILLER_24_307 ();
 decap_12 FILLER_24_309 ();
 decap_12 FILLER_24_321 ();
 decap_12 FILLER_24_333 ();
 decap_12 FILLER_24_345 ();
 fill_4 FILLER_24_357 ();
 fill_2 FILLER_24_361 ();
 fill_1 FILLER_24_363 ();
 decap_12 FILLER_24_365 ();
 decap_12 FILLER_24_377 ();
 decap_12 FILLER_24_389 ();
 decap_12 FILLER_24_401 ();
 fill_4 FILLER_24_413 ();
 fill_2 FILLER_24_417 ();
 fill_1 FILLER_24_419 ();
 decap_12 FILLER_24_421 ();
 decap_12 FILLER_24_433 ();
 decap_12 FILLER_24_445 ();
 decap_12 FILLER_24_457 ();
 fill_4 FILLER_24_469 ();
 fill_2 FILLER_24_473 ();
 fill_1 FILLER_24_475 ();
 decap_12 FILLER_24_477 ();
 decap_12 FILLER_24_489 ();
 decap_12 FILLER_24_501 ();
 decap_12 FILLER_24_513 ();
 fill_4 FILLER_24_525 ();
 fill_2 FILLER_24_529 ();
 fill_1 FILLER_24_531 ();
 decap_12 FILLER_24_533 ();
 decap_12 FILLER_24_545 ();
 decap_12 FILLER_24_557 ();
 decap_12 FILLER_24_569 ();
 fill_4 FILLER_24_581 ();
 fill_2 FILLER_24_585 ();
 fill_1 FILLER_24_587 ();
 decap_12 FILLER_24_589 ();
 decap_12 FILLER_24_601 ();
 decap_12 FILLER_24_613 ();
 decap_12 FILLER_25_3 ();
 decap_12 FILLER_25_15 ();
 decap_12 FILLER_25_27 ();
 decap_12 FILLER_25_39 ();
 fill_4 FILLER_25_51 ();
 fill_1 FILLER_25_55 ();
 decap_12 FILLER_25_57 ();
 decap_12 FILLER_25_69 ();
 decap_12 FILLER_25_81 ();
 decap_12 FILLER_25_93 ();
 fill_4 FILLER_25_105 ();
 fill_2 FILLER_25_109 ();
 fill_1 FILLER_25_111 ();
 decap_12 FILLER_25_113 ();
 decap_12 FILLER_25_125 ();
 decap_12 FILLER_25_137 ();
 decap_12 FILLER_25_149 ();
 fill_4 FILLER_25_161 ();
 fill_2 FILLER_25_165 ();
 fill_1 FILLER_25_167 ();
 decap_12 FILLER_25_169 ();
 decap_12 FILLER_25_181 ();
 decap_12 FILLER_25_193 ();
 decap_12 FILLER_25_205 ();
 fill_4 FILLER_25_217 ();
 fill_2 FILLER_25_221 ();
 fill_1 FILLER_25_223 ();
 decap_12 FILLER_25_225 ();
 decap_12 FILLER_25_237 ();
 decap_12 FILLER_25_249 ();
 decap_12 FILLER_25_261 ();
 fill_4 FILLER_25_273 ();
 fill_2 FILLER_25_277 ();
 fill_1 FILLER_25_279 ();
 decap_12 FILLER_25_281 ();
 decap_12 FILLER_25_293 ();
 decap_12 FILLER_25_305 ();
 decap_12 FILLER_25_317 ();
 fill_4 FILLER_25_329 ();
 fill_2 FILLER_25_333 ();
 fill_1 FILLER_25_335 ();
 decap_12 FILLER_25_337 ();
 decap_12 FILLER_25_349 ();
 decap_12 FILLER_25_361 ();
 decap_12 FILLER_25_373 ();
 fill_4 FILLER_25_385 ();
 fill_2 FILLER_25_389 ();
 fill_1 FILLER_25_391 ();
 decap_12 FILLER_25_393 ();
 decap_12 FILLER_25_405 ();
 decap_12 FILLER_25_417 ();
 decap_12 FILLER_25_429 ();
 fill_4 FILLER_25_441 ();
 fill_2 FILLER_25_445 ();
 fill_1 FILLER_25_447 ();
 decap_12 FILLER_25_449 ();
 decap_12 FILLER_25_461 ();
 decap_12 FILLER_25_473 ();
 decap_12 FILLER_25_485 ();
 fill_4 FILLER_25_497 ();
 fill_2 FILLER_25_501 ();
 fill_1 FILLER_25_503 ();
 decap_12 FILLER_25_505 ();
 decap_12 FILLER_25_517 ();
 decap_12 FILLER_25_529 ();
 decap_12 FILLER_25_541 ();
 fill_4 FILLER_25_553 ();
 fill_2 FILLER_25_557 ();
 fill_1 FILLER_25_559 ();
 decap_12 FILLER_25_561 ();
 decap_12 FILLER_25_573 ();
 decap_12 FILLER_25_585 ();
 decap_12 FILLER_25_597 ();
 fill_4 FILLER_25_609 ();
 fill_2 FILLER_25_613 ();
 fill_1 FILLER_25_615 ();
 fill_8 FILLER_25_617 ();
 decap_12 FILLER_26_3 ();
 decap_12 FILLER_26_15 ();
 fill_1 FILLER_26_27 ();
 decap_12 FILLER_26_29 ();
 decap_12 FILLER_26_41 ();
 decap_12 FILLER_26_53 ();
 decap_12 FILLER_26_65 ();
 fill_4 FILLER_26_77 ();
 fill_2 FILLER_26_81 ();
 fill_1 FILLER_26_83 ();
 decap_12 FILLER_26_85 ();
 decap_12 FILLER_26_97 ();
 decap_12 FILLER_26_109 ();
 decap_12 FILLER_26_121 ();
 fill_4 FILLER_26_133 ();
 fill_2 FILLER_26_137 ();
 fill_1 FILLER_26_139 ();
 decap_12 FILLER_26_141 ();
 decap_12 FILLER_26_153 ();
 decap_12 FILLER_26_165 ();
 decap_12 FILLER_26_177 ();
 fill_4 FILLER_26_189 ();
 fill_2 FILLER_26_193 ();
 fill_1 FILLER_26_195 ();
 decap_12 FILLER_26_197 ();
 decap_12 FILLER_26_209 ();
 decap_12 FILLER_26_221 ();
 decap_12 FILLER_26_233 ();
 fill_4 FILLER_26_245 ();
 fill_2 FILLER_26_249 ();
 fill_1 FILLER_26_251 ();
 decap_12 FILLER_26_253 ();
 decap_12 FILLER_26_265 ();
 decap_12 FILLER_26_277 ();
 decap_12 FILLER_26_289 ();
 fill_4 FILLER_26_301 ();
 fill_2 FILLER_26_305 ();
 fill_1 FILLER_26_307 ();
 decap_12 FILLER_26_309 ();
 decap_12 FILLER_26_321 ();
 decap_12 FILLER_26_333 ();
 decap_12 FILLER_26_345 ();
 fill_4 FILLER_26_357 ();
 fill_2 FILLER_26_361 ();
 fill_1 FILLER_26_363 ();
 decap_12 FILLER_26_365 ();
 decap_12 FILLER_26_377 ();
 decap_12 FILLER_26_389 ();
 decap_12 FILLER_26_401 ();
 fill_4 FILLER_26_413 ();
 fill_2 FILLER_26_417 ();
 fill_1 FILLER_26_419 ();
 decap_12 FILLER_26_421 ();
 decap_12 FILLER_26_433 ();
 decap_12 FILLER_26_445 ();
 decap_12 FILLER_26_457 ();
 fill_4 FILLER_26_469 ();
 fill_2 FILLER_26_473 ();
 fill_1 FILLER_26_475 ();
 decap_12 FILLER_26_477 ();
 decap_12 FILLER_26_489 ();
 decap_12 FILLER_26_501 ();
 decap_12 FILLER_26_513 ();
 fill_4 FILLER_26_525 ();
 fill_2 FILLER_26_529 ();
 fill_1 FILLER_26_531 ();
 decap_12 FILLER_26_533 ();
 decap_12 FILLER_26_545 ();
 decap_12 FILLER_26_557 ();
 decap_12 FILLER_26_569 ();
 fill_4 FILLER_26_581 ();
 fill_2 FILLER_26_585 ();
 fill_1 FILLER_26_587 ();
 decap_12 FILLER_26_589 ();
 decap_12 FILLER_26_601 ();
 decap_12 FILLER_26_613 ();
 decap_12 FILLER_27_3 ();
 decap_12 FILLER_27_15 ();
 decap_12 FILLER_27_27 ();
 decap_12 FILLER_27_39 ();
 fill_4 FILLER_27_51 ();
 fill_1 FILLER_27_55 ();
 decap_12 FILLER_27_57 ();
 decap_12 FILLER_27_69 ();
 decap_12 FILLER_27_81 ();
 decap_12 FILLER_27_93 ();
 fill_4 FILLER_27_105 ();
 fill_2 FILLER_27_109 ();
 fill_1 FILLER_27_111 ();
 decap_12 FILLER_27_113 ();
 decap_12 FILLER_27_125 ();
 decap_12 FILLER_27_137 ();
 decap_12 FILLER_27_149 ();
 fill_4 FILLER_27_161 ();
 fill_2 FILLER_27_165 ();
 fill_1 FILLER_27_167 ();
 decap_12 FILLER_27_169 ();
 decap_12 FILLER_27_181 ();
 decap_12 FILLER_27_193 ();
 decap_12 FILLER_27_205 ();
 fill_4 FILLER_27_217 ();
 fill_2 FILLER_27_221 ();
 fill_1 FILLER_27_223 ();
 decap_12 FILLER_27_225 ();
 decap_12 FILLER_27_237 ();
 decap_12 FILLER_27_249 ();
 decap_12 FILLER_27_261 ();
 fill_4 FILLER_27_273 ();
 fill_2 FILLER_27_277 ();
 fill_1 FILLER_27_279 ();
 decap_12 FILLER_27_281 ();
 decap_12 FILLER_27_293 ();
 decap_12 FILLER_27_305 ();
 decap_12 FILLER_27_317 ();
 fill_4 FILLER_27_329 ();
 fill_2 FILLER_27_333 ();
 fill_1 FILLER_27_335 ();
 decap_12 FILLER_27_337 ();
 decap_12 FILLER_27_349 ();
 decap_12 FILLER_27_361 ();
 decap_12 FILLER_27_373 ();
 fill_4 FILLER_27_385 ();
 fill_2 FILLER_27_389 ();
 fill_1 FILLER_27_391 ();
 decap_12 FILLER_27_393 ();
 decap_12 FILLER_27_405 ();
 decap_12 FILLER_27_417 ();
 decap_12 FILLER_27_429 ();
 fill_4 FILLER_27_441 ();
 fill_2 FILLER_27_445 ();
 fill_1 FILLER_27_447 ();
 decap_12 FILLER_27_449 ();
 decap_12 FILLER_27_461 ();
 decap_12 FILLER_27_473 ();
 decap_12 FILLER_27_485 ();
 fill_4 FILLER_27_497 ();
 fill_2 FILLER_27_501 ();
 fill_1 FILLER_27_503 ();
 decap_12 FILLER_27_505 ();
 decap_12 FILLER_27_517 ();
 decap_12 FILLER_27_529 ();
 decap_12 FILLER_27_541 ();
 fill_4 FILLER_27_553 ();
 fill_2 FILLER_27_557 ();
 fill_1 FILLER_27_559 ();
 decap_12 FILLER_27_561 ();
 decap_12 FILLER_27_573 ();
 decap_12 FILLER_27_585 ();
 decap_12 FILLER_27_597 ();
 fill_4 FILLER_27_609 ();
 fill_2 FILLER_27_613 ();
 fill_1 FILLER_27_615 ();
 fill_8 FILLER_27_617 ();
 decap_12 FILLER_28_3 ();
 decap_12 FILLER_28_15 ();
 fill_1 FILLER_28_27 ();
 decap_12 FILLER_28_29 ();
 decap_12 FILLER_28_41 ();
 decap_12 FILLER_28_53 ();
 decap_12 FILLER_28_65 ();
 fill_4 FILLER_28_77 ();
 fill_2 FILLER_28_81 ();
 fill_1 FILLER_28_83 ();
 decap_12 FILLER_28_85 ();
 decap_12 FILLER_28_97 ();
 decap_12 FILLER_28_109 ();
 decap_12 FILLER_28_121 ();
 fill_4 FILLER_28_133 ();
 fill_2 FILLER_28_137 ();
 fill_1 FILLER_28_139 ();
 decap_12 FILLER_28_141 ();
 decap_12 FILLER_28_153 ();
 decap_12 FILLER_28_165 ();
 decap_12 FILLER_28_177 ();
 fill_4 FILLER_28_189 ();
 fill_2 FILLER_28_193 ();
 fill_1 FILLER_28_195 ();
 decap_12 FILLER_28_197 ();
 decap_12 FILLER_28_209 ();
 decap_12 FILLER_28_221 ();
 decap_12 FILLER_28_233 ();
 fill_4 FILLER_28_245 ();
 fill_2 FILLER_28_249 ();
 fill_1 FILLER_28_251 ();
 decap_12 FILLER_28_253 ();
 decap_12 FILLER_28_265 ();
 decap_12 FILLER_28_277 ();
 decap_12 FILLER_28_289 ();
 fill_4 FILLER_28_301 ();
 fill_2 FILLER_28_305 ();
 fill_1 FILLER_28_307 ();
 decap_12 FILLER_28_309 ();
 decap_12 FILLER_28_321 ();
 decap_12 FILLER_28_333 ();
 decap_12 FILLER_28_345 ();
 fill_4 FILLER_28_357 ();
 fill_2 FILLER_28_361 ();
 fill_1 FILLER_28_363 ();
 decap_12 FILLER_28_365 ();
 decap_12 FILLER_28_377 ();
 decap_12 FILLER_28_389 ();
 decap_12 FILLER_28_401 ();
 fill_4 FILLER_28_413 ();
 fill_2 FILLER_28_417 ();
 fill_1 FILLER_28_419 ();
 decap_12 FILLER_28_421 ();
 decap_12 FILLER_28_433 ();
 decap_12 FILLER_28_445 ();
 decap_12 FILLER_28_457 ();
 fill_4 FILLER_28_469 ();
 fill_2 FILLER_28_473 ();
 fill_1 FILLER_28_475 ();
 decap_12 FILLER_28_477 ();
 decap_12 FILLER_28_489 ();
 decap_12 FILLER_28_501 ();
 decap_12 FILLER_28_513 ();
 fill_4 FILLER_28_525 ();
 fill_2 FILLER_28_529 ();
 fill_1 FILLER_28_531 ();
 decap_12 FILLER_28_533 ();
 decap_12 FILLER_28_545 ();
 decap_12 FILLER_28_557 ();
 decap_12 FILLER_28_569 ();
 fill_4 FILLER_28_581 ();
 fill_2 FILLER_28_585 ();
 fill_1 FILLER_28_587 ();
 decap_12 FILLER_28_589 ();
 decap_12 FILLER_28_601 ();
 decap_12 FILLER_28_613 ();
 decap_12 FILLER_29_3 ();
 decap_12 FILLER_29_15 ();
 decap_12 FILLER_29_27 ();
 decap_12 FILLER_29_39 ();
 fill_4 FILLER_29_51 ();
 fill_1 FILLER_29_55 ();
 decap_12 FILLER_29_57 ();
 decap_12 FILLER_29_69 ();
 decap_12 FILLER_29_81 ();
 decap_12 FILLER_29_93 ();
 fill_4 FILLER_29_105 ();
 fill_2 FILLER_29_109 ();
 fill_1 FILLER_29_111 ();
 decap_12 FILLER_29_113 ();
 decap_12 FILLER_29_125 ();
 decap_12 FILLER_29_137 ();
 decap_12 FILLER_29_149 ();
 fill_4 FILLER_29_161 ();
 fill_2 FILLER_29_165 ();
 fill_1 FILLER_29_167 ();
 decap_12 FILLER_29_169 ();
 decap_12 FILLER_29_181 ();
 decap_12 FILLER_29_193 ();
 decap_12 FILLER_29_205 ();
 fill_4 FILLER_29_217 ();
 fill_2 FILLER_29_221 ();
 fill_1 FILLER_29_223 ();
 decap_12 FILLER_29_225 ();
 decap_12 FILLER_29_237 ();
 decap_12 FILLER_29_249 ();
 decap_12 FILLER_29_261 ();
 fill_4 FILLER_29_273 ();
 fill_2 FILLER_29_277 ();
 fill_1 FILLER_29_279 ();
 decap_12 FILLER_29_281 ();
 decap_12 FILLER_29_293 ();
 decap_12 FILLER_29_305 ();
 decap_12 FILLER_29_317 ();
 fill_4 FILLER_29_329 ();
 fill_2 FILLER_29_333 ();
 fill_1 FILLER_29_335 ();
 decap_12 FILLER_29_337 ();
 decap_12 FILLER_29_349 ();
 decap_12 FILLER_29_361 ();
 decap_12 FILLER_29_373 ();
 fill_4 FILLER_29_385 ();
 fill_2 FILLER_29_389 ();
 fill_1 FILLER_29_391 ();
 decap_12 FILLER_29_393 ();
 decap_12 FILLER_29_405 ();
 decap_12 FILLER_29_417 ();
 decap_12 FILLER_29_429 ();
 fill_4 FILLER_29_441 ();
 fill_2 FILLER_29_445 ();
 fill_1 FILLER_29_447 ();
 decap_12 FILLER_29_449 ();
 decap_12 FILLER_29_461 ();
 decap_12 FILLER_29_473 ();
 decap_12 FILLER_29_485 ();
 fill_4 FILLER_29_497 ();
 fill_2 FILLER_29_501 ();
 fill_1 FILLER_29_503 ();
 decap_12 FILLER_29_505 ();
 decap_12 FILLER_29_517 ();
 decap_12 FILLER_29_529 ();
 decap_12 FILLER_29_541 ();
 fill_4 FILLER_29_553 ();
 fill_2 FILLER_29_557 ();
 fill_1 FILLER_29_559 ();
 decap_12 FILLER_29_561 ();
 decap_12 FILLER_29_573 ();
 decap_12 FILLER_29_585 ();
 decap_12 FILLER_29_597 ();
 fill_4 FILLER_29_609 ();
 fill_2 FILLER_29_613 ();
 fill_1 FILLER_29_615 ();
 fill_8 FILLER_29_617 ();
 decap_12 FILLER_30_3 ();
 decap_12 FILLER_30_15 ();
 fill_1 FILLER_30_27 ();
 decap_12 FILLER_30_29 ();
 decap_12 FILLER_30_41 ();
 decap_12 FILLER_30_53 ();
 decap_12 FILLER_30_65 ();
 fill_4 FILLER_30_77 ();
 fill_2 FILLER_30_81 ();
 fill_1 FILLER_30_83 ();
 decap_12 FILLER_30_85 ();
 decap_12 FILLER_30_97 ();
 decap_12 FILLER_30_109 ();
 decap_12 FILLER_30_121 ();
 fill_4 FILLER_30_133 ();
 fill_2 FILLER_30_137 ();
 fill_1 FILLER_30_139 ();
 decap_12 FILLER_30_141 ();
 decap_12 FILLER_30_153 ();
 decap_12 FILLER_30_165 ();
 decap_12 FILLER_30_177 ();
 fill_4 FILLER_30_189 ();
 fill_2 FILLER_30_193 ();
 fill_1 FILLER_30_195 ();
 decap_12 FILLER_30_197 ();
 decap_12 FILLER_30_209 ();
 decap_12 FILLER_30_221 ();
 decap_12 FILLER_30_233 ();
 fill_4 FILLER_30_245 ();
 fill_2 FILLER_30_249 ();
 fill_1 FILLER_30_251 ();
 decap_12 FILLER_30_253 ();
 decap_12 FILLER_30_265 ();
 decap_12 FILLER_30_277 ();
 decap_12 FILLER_30_289 ();
 fill_4 FILLER_30_301 ();
 fill_2 FILLER_30_305 ();
 fill_1 FILLER_30_307 ();
 decap_12 FILLER_30_309 ();
 decap_12 FILLER_30_321 ();
 decap_12 FILLER_30_333 ();
 decap_12 FILLER_30_345 ();
 fill_4 FILLER_30_357 ();
 fill_2 FILLER_30_361 ();
 fill_1 FILLER_30_363 ();
 decap_12 FILLER_30_365 ();
 decap_12 FILLER_30_377 ();
 decap_12 FILLER_30_389 ();
 decap_12 FILLER_30_401 ();
 fill_4 FILLER_30_413 ();
 fill_2 FILLER_30_417 ();
 fill_1 FILLER_30_419 ();
 decap_12 FILLER_30_421 ();
 decap_12 FILLER_30_433 ();
 decap_12 FILLER_30_445 ();
 decap_12 FILLER_30_457 ();
 fill_4 FILLER_30_469 ();
 fill_2 FILLER_30_473 ();
 fill_1 FILLER_30_475 ();
 decap_12 FILLER_30_477 ();
 decap_12 FILLER_30_489 ();
 decap_12 FILLER_30_501 ();
 decap_12 FILLER_30_513 ();
 fill_4 FILLER_30_525 ();
 fill_2 FILLER_30_529 ();
 fill_1 FILLER_30_531 ();
 decap_12 FILLER_30_533 ();
 decap_12 FILLER_30_545 ();
 decap_12 FILLER_30_557 ();
 decap_12 FILLER_30_569 ();
 fill_4 FILLER_30_581 ();
 fill_2 FILLER_30_585 ();
 fill_1 FILLER_30_587 ();
 decap_12 FILLER_30_589 ();
 decap_12 FILLER_30_601 ();
 decap_12 FILLER_30_613 ();
 decap_12 FILLER_31_3 ();
 decap_12 FILLER_31_15 ();
 decap_12 FILLER_31_27 ();
 decap_12 FILLER_31_39 ();
 fill_4 FILLER_31_51 ();
 fill_1 FILLER_31_55 ();
 decap_12 FILLER_31_57 ();
 decap_12 FILLER_31_69 ();
 decap_12 FILLER_31_81 ();
 decap_12 FILLER_31_93 ();
 fill_4 FILLER_31_105 ();
 fill_2 FILLER_31_109 ();
 fill_1 FILLER_31_111 ();
 decap_12 FILLER_31_113 ();
 decap_12 FILLER_31_125 ();
 decap_12 FILLER_31_137 ();
 decap_12 FILLER_31_149 ();
 fill_4 FILLER_31_161 ();
 fill_2 FILLER_31_165 ();
 fill_1 FILLER_31_167 ();
 decap_12 FILLER_31_169 ();
 decap_12 FILLER_31_181 ();
 decap_12 FILLER_31_193 ();
 decap_12 FILLER_31_205 ();
 fill_4 FILLER_31_217 ();
 fill_2 FILLER_31_221 ();
 fill_1 FILLER_31_223 ();
 decap_12 FILLER_31_225 ();
 decap_12 FILLER_31_237 ();
 decap_12 FILLER_31_249 ();
 decap_12 FILLER_31_261 ();
 fill_4 FILLER_31_273 ();
 fill_2 FILLER_31_277 ();
 fill_1 FILLER_31_279 ();
 decap_12 FILLER_31_281 ();
 decap_12 FILLER_31_293 ();
 decap_12 FILLER_31_305 ();
 decap_12 FILLER_31_317 ();
 fill_4 FILLER_31_329 ();
 fill_2 FILLER_31_333 ();
 fill_1 FILLER_31_335 ();
 decap_12 FILLER_31_337 ();
 decap_12 FILLER_31_349 ();
 decap_12 FILLER_31_361 ();
 decap_12 FILLER_31_373 ();
 fill_4 FILLER_31_385 ();
 fill_2 FILLER_31_389 ();
 fill_1 FILLER_31_391 ();
 decap_12 FILLER_31_393 ();
 decap_12 FILLER_31_405 ();
 decap_12 FILLER_31_417 ();
 decap_12 FILLER_31_429 ();
 fill_4 FILLER_31_441 ();
 fill_2 FILLER_31_445 ();
 fill_1 FILLER_31_447 ();
 decap_12 FILLER_31_449 ();
 decap_12 FILLER_31_461 ();
 decap_12 FILLER_31_473 ();
 decap_12 FILLER_31_485 ();
 fill_4 FILLER_31_497 ();
 fill_2 FILLER_31_501 ();
 fill_1 FILLER_31_503 ();
 decap_12 FILLER_31_505 ();
 decap_12 FILLER_31_517 ();
 decap_12 FILLER_31_529 ();
 decap_12 FILLER_31_541 ();
 fill_4 FILLER_31_553 ();
 fill_2 FILLER_31_557 ();
 fill_1 FILLER_31_559 ();
 decap_12 FILLER_31_561 ();
 decap_12 FILLER_31_573 ();
 decap_12 FILLER_31_585 ();
 decap_12 FILLER_31_597 ();
 fill_4 FILLER_31_609 ();
 fill_2 FILLER_31_613 ();
 fill_1 FILLER_31_615 ();
 fill_8 FILLER_31_617 ();
 decap_12 FILLER_32_3 ();
 decap_12 FILLER_32_15 ();
 fill_1 FILLER_32_27 ();
 decap_12 FILLER_32_29 ();
 decap_12 FILLER_32_41 ();
 decap_12 FILLER_32_53 ();
 decap_12 FILLER_32_65 ();
 fill_4 FILLER_32_77 ();
 fill_2 FILLER_32_81 ();
 fill_1 FILLER_32_83 ();
 decap_12 FILLER_32_85 ();
 decap_12 FILLER_32_97 ();
 decap_12 FILLER_32_109 ();
 decap_12 FILLER_32_121 ();
 fill_4 FILLER_32_133 ();
 fill_2 FILLER_32_137 ();
 fill_1 FILLER_32_139 ();
 decap_12 FILLER_32_141 ();
 decap_12 FILLER_32_153 ();
 decap_12 FILLER_32_165 ();
 decap_12 FILLER_32_177 ();
 fill_4 FILLER_32_189 ();
 fill_2 FILLER_32_193 ();
 fill_1 FILLER_32_195 ();
 decap_12 FILLER_32_197 ();
 decap_12 FILLER_32_209 ();
 decap_12 FILLER_32_221 ();
 decap_12 FILLER_32_233 ();
 fill_4 FILLER_32_245 ();
 fill_2 FILLER_32_249 ();
 fill_1 FILLER_32_251 ();
 decap_12 FILLER_32_253 ();
 decap_12 FILLER_32_265 ();
 decap_12 FILLER_32_277 ();
 decap_12 FILLER_32_289 ();
 fill_4 FILLER_32_301 ();
 fill_2 FILLER_32_305 ();
 fill_1 FILLER_32_307 ();
 decap_12 FILLER_32_309 ();
 decap_12 FILLER_32_321 ();
 decap_12 FILLER_32_333 ();
 decap_12 FILLER_32_345 ();
 fill_4 FILLER_32_357 ();
 fill_2 FILLER_32_361 ();
 fill_1 FILLER_32_363 ();
 decap_12 FILLER_32_365 ();
 decap_12 FILLER_32_377 ();
 decap_12 FILLER_32_389 ();
 decap_12 FILLER_32_401 ();
 fill_4 FILLER_32_413 ();
 fill_2 FILLER_32_417 ();
 fill_1 FILLER_32_419 ();
 decap_12 FILLER_32_421 ();
 decap_12 FILLER_32_433 ();
 decap_12 FILLER_32_445 ();
 decap_12 FILLER_32_457 ();
 fill_4 FILLER_32_469 ();
 fill_2 FILLER_32_473 ();
 fill_1 FILLER_32_475 ();
 decap_12 FILLER_32_477 ();
 decap_12 FILLER_32_489 ();
 decap_12 FILLER_32_501 ();
 decap_12 FILLER_32_513 ();
 fill_4 FILLER_32_525 ();
 fill_2 FILLER_32_529 ();
 fill_1 FILLER_32_531 ();
 decap_12 FILLER_32_533 ();
 decap_12 FILLER_32_545 ();
 decap_12 FILLER_32_557 ();
 decap_12 FILLER_32_569 ();
 fill_4 FILLER_32_581 ();
 fill_2 FILLER_32_585 ();
 fill_1 FILLER_32_587 ();
 decap_12 FILLER_32_589 ();
 decap_12 FILLER_32_601 ();
 decap_12 FILLER_32_613 ();
 decap_12 FILLER_33_3 ();
 decap_12 FILLER_33_15 ();
 decap_12 FILLER_33_27 ();
 decap_12 FILLER_33_39 ();
 fill_4 FILLER_33_51 ();
 fill_1 FILLER_33_55 ();
 decap_12 FILLER_33_57 ();
 decap_12 FILLER_33_69 ();
 decap_12 FILLER_33_81 ();
 decap_12 FILLER_33_93 ();
 fill_4 FILLER_33_105 ();
 fill_2 FILLER_33_109 ();
 fill_1 FILLER_33_111 ();
 decap_12 FILLER_33_113 ();
 decap_12 FILLER_33_125 ();
 decap_12 FILLER_33_137 ();
 decap_12 FILLER_33_149 ();
 fill_4 FILLER_33_161 ();
 fill_2 FILLER_33_165 ();
 fill_1 FILLER_33_167 ();
 decap_12 FILLER_33_169 ();
 decap_12 FILLER_33_181 ();
 decap_12 FILLER_33_193 ();
 decap_12 FILLER_33_205 ();
 fill_4 FILLER_33_217 ();
 fill_2 FILLER_33_221 ();
 fill_1 FILLER_33_223 ();
 decap_12 FILLER_33_225 ();
 decap_12 FILLER_33_237 ();
 decap_12 FILLER_33_249 ();
 decap_12 FILLER_33_261 ();
 fill_4 FILLER_33_273 ();
 fill_2 FILLER_33_277 ();
 fill_1 FILLER_33_279 ();
 decap_12 FILLER_33_281 ();
 decap_12 FILLER_33_293 ();
 decap_12 FILLER_33_305 ();
 decap_12 FILLER_33_317 ();
 fill_4 FILLER_33_329 ();
 fill_2 FILLER_33_333 ();
 fill_1 FILLER_33_335 ();
 decap_12 FILLER_33_337 ();
 decap_12 FILLER_33_349 ();
 decap_12 FILLER_33_361 ();
 decap_12 FILLER_33_373 ();
 fill_4 FILLER_33_385 ();
 fill_2 FILLER_33_389 ();
 fill_1 FILLER_33_391 ();
 decap_12 FILLER_33_393 ();
 decap_12 FILLER_33_405 ();
 decap_12 FILLER_33_417 ();
 decap_12 FILLER_33_429 ();
 fill_4 FILLER_33_441 ();
 fill_2 FILLER_33_445 ();
 fill_1 FILLER_33_447 ();
 decap_12 FILLER_33_449 ();
 decap_12 FILLER_33_461 ();
 decap_12 FILLER_33_473 ();
 decap_12 FILLER_33_485 ();
 fill_4 FILLER_33_497 ();
 fill_2 FILLER_33_501 ();
 fill_1 FILLER_33_503 ();
 decap_12 FILLER_33_505 ();
 decap_12 FILLER_33_517 ();
 decap_12 FILLER_33_529 ();
 decap_12 FILLER_33_541 ();
 fill_4 FILLER_33_553 ();
 fill_2 FILLER_33_557 ();
 fill_1 FILLER_33_559 ();
 decap_12 FILLER_33_561 ();
 decap_12 FILLER_33_573 ();
 decap_12 FILLER_33_585 ();
 decap_12 FILLER_33_597 ();
 fill_4 FILLER_33_609 ();
 fill_2 FILLER_33_613 ();
 fill_1 FILLER_33_615 ();
 fill_8 FILLER_33_617 ();
 decap_12 FILLER_34_3 ();
 decap_12 FILLER_34_15 ();
 fill_1 FILLER_34_27 ();
 decap_12 FILLER_34_29 ();
 decap_12 FILLER_34_41 ();
 decap_12 FILLER_34_53 ();
 decap_12 FILLER_34_65 ();
 fill_4 FILLER_34_77 ();
 fill_2 FILLER_34_81 ();
 fill_1 FILLER_34_83 ();
 decap_12 FILLER_34_85 ();
 decap_12 FILLER_34_97 ();
 decap_12 FILLER_34_109 ();
 decap_12 FILLER_34_121 ();
 fill_4 FILLER_34_133 ();
 fill_2 FILLER_34_137 ();
 fill_1 FILLER_34_139 ();
 decap_12 FILLER_34_141 ();
 decap_12 FILLER_34_153 ();
 decap_12 FILLER_34_165 ();
 decap_12 FILLER_34_177 ();
 fill_4 FILLER_34_189 ();
 fill_2 FILLER_34_193 ();
 fill_1 FILLER_34_195 ();
 decap_12 FILLER_34_197 ();
 decap_12 FILLER_34_209 ();
 decap_12 FILLER_34_221 ();
 decap_12 FILLER_34_233 ();
 fill_4 FILLER_34_245 ();
 fill_2 FILLER_34_249 ();
 fill_1 FILLER_34_251 ();
 decap_12 FILLER_34_253 ();
 decap_12 FILLER_34_265 ();
 decap_12 FILLER_34_277 ();
 decap_12 FILLER_34_289 ();
 fill_4 FILLER_34_301 ();
 fill_2 FILLER_34_305 ();
 fill_1 FILLER_34_307 ();
 decap_12 FILLER_34_309 ();
 decap_12 FILLER_34_321 ();
 decap_12 FILLER_34_333 ();
 decap_12 FILLER_34_345 ();
 fill_4 FILLER_34_357 ();
 fill_2 FILLER_34_361 ();
 fill_1 FILLER_34_363 ();
 decap_12 FILLER_34_365 ();
 decap_12 FILLER_34_377 ();
 decap_12 FILLER_34_389 ();
 decap_12 FILLER_34_401 ();
 fill_4 FILLER_34_413 ();
 fill_2 FILLER_34_417 ();
 fill_1 FILLER_34_419 ();
 decap_12 FILLER_34_421 ();
 decap_12 FILLER_34_433 ();
 decap_12 FILLER_34_445 ();
 decap_12 FILLER_34_457 ();
 fill_4 FILLER_34_469 ();
 fill_2 FILLER_34_473 ();
 fill_1 FILLER_34_475 ();
 decap_12 FILLER_34_477 ();
 decap_12 FILLER_34_489 ();
 decap_12 FILLER_34_501 ();
 decap_12 FILLER_34_513 ();
 fill_4 FILLER_34_525 ();
 fill_2 FILLER_34_529 ();
 fill_1 FILLER_34_531 ();
 decap_12 FILLER_34_533 ();
 decap_12 FILLER_34_545 ();
 decap_12 FILLER_34_557 ();
 decap_12 FILLER_34_569 ();
 fill_4 FILLER_34_581 ();
 fill_2 FILLER_34_585 ();
 fill_1 FILLER_34_587 ();
 decap_12 FILLER_34_589 ();
 decap_12 FILLER_34_601 ();
 decap_12 FILLER_34_613 ();
 decap_12 FILLER_35_3 ();
 decap_12 FILLER_35_15 ();
 decap_12 FILLER_35_27 ();
 decap_12 FILLER_35_39 ();
 fill_4 FILLER_35_51 ();
 fill_1 FILLER_35_55 ();
 decap_12 FILLER_35_57 ();
 decap_12 FILLER_35_69 ();
 decap_12 FILLER_35_81 ();
 decap_12 FILLER_35_93 ();
 fill_4 FILLER_35_105 ();
 fill_2 FILLER_35_109 ();
 fill_1 FILLER_35_111 ();
 decap_12 FILLER_35_113 ();
 decap_12 FILLER_35_125 ();
 decap_12 FILLER_35_137 ();
 decap_12 FILLER_35_149 ();
 fill_4 FILLER_35_161 ();
 fill_2 FILLER_35_165 ();
 fill_1 FILLER_35_167 ();
 decap_12 FILLER_35_169 ();
 decap_12 FILLER_35_181 ();
 decap_12 FILLER_35_193 ();
 decap_12 FILLER_35_205 ();
 fill_4 FILLER_35_217 ();
 fill_2 FILLER_35_221 ();
 fill_1 FILLER_35_223 ();
 decap_12 FILLER_35_225 ();
 decap_12 FILLER_35_237 ();
 decap_12 FILLER_35_249 ();
 decap_12 FILLER_35_261 ();
 fill_4 FILLER_35_273 ();
 fill_2 FILLER_35_277 ();
 fill_1 FILLER_35_279 ();
 decap_12 FILLER_35_281 ();
 decap_12 FILLER_35_293 ();
 decap_12 FILLER_35_305 ();
 decap_12 FILLER_35_317 ();
 fill_4 FILLER_35_329 ();
 fill_2 FILLER_35_333 ();
 fill_1 FILLER_35_335 ();
 decap_12 FILLER_35_337 ();
 decap_12 FILLER_35_349 ();
 decap_12 FILLER_35_361 ();
 decap_12 FILLER_35_373 ();
 fill_4 FILLER_35_385 ();
 fill_2 FILLER_35_389 ();
 fill_1 FILLER_35_391 ();
 decap_12 FILLER_35_393 ();
 decap_12 FILLER_35_405 ();
 decap_12 FILLER_35_417 ();
 decap_12 FILLER_35_429 ();
 fill_4 FILLER_35_441 ();
 fill_2 FILLER_35_445 ();
 fill_1 FILLER_35_447 ();
 decap_12 FILLER_35_449 ();
 decap_12 FILLER_35_461 ();
 decap_12 FILLER_35_473 ();
 decap_12 FILLER_35_485 ();
 fill_4 FILLER_35_497 ();
 fill_2 FILLER_35_501 ();
 fill_1 FILLER_35_503 ();
 decap_12 FILLER_35_505 ();
 decap_12 FILLER_35_517 ();
 decap_12 FILLER_35_529 ();
 decap_12 FILLER_35_541 ();
 fill_4 FILLER_35_553 ();
 fill_2 FILLER_35_557 ();
 fill_1 FILLER_35_559 ();
 decap_12 FILLER_35_561 ();
 decap_12 FILLER_35_573 ();
 decap_12 FILLER_35_585 ();
 decap_12 FILLER_35_597 ();
 fill_4 FILLER_35_609 ();
 fill_2 FILLER_35_613 ();
 fill_1 FILLER_35_615 ();
 fill_8 FILLER_35_617 ();
 decap_12 FILLER_36_3 ();
 decap_12 FILLER_36_15 ();
 fill_1 FILLER_36_27 ();
 decap_12 FILLER_36_29 ();
 decap_12 FILLER_36_41 ();
 decap_12 FILLER_36_53 ();
 decap_12 FILLER_36_65 ();
 fill_4 FILLER_36_77 ();
 fill_2 FILLER_36_81 ();
 fill_1 FILLER_36_83 ();
 decap_12 FILLER_36_85 ();
 decap_12 FILLER_36_97 ();
 decap_12 FILLER_36_109 ();
 decap_12 FILLER_36_121 ();
 fill_4 FILLER_36_133 ();
 fill_2 FILLER_36_137 ();
 fill_1 FILLER_36_139 ();
 decap_12 FILLER_36_141 ();
 decap_12 FILLER_36_153 ();
 decap_12 FILLER_36_165 ();
 decap_12 FILLER_36_177 ();
 fill_4 FILLER_36_189 ();
 fill_2 FILLER_36_193 ();
 fill_1 FILLER_36_195 ();
 decap_12 FILLER_36_197 ();
 decap_12 FILLER_36_209 ();
 decap_12 FILLER_36_221 ();
 decap_12 FILLER_36_233 ();
 fill_4 FILLER_36_245 ();
 fill_2 FILLER_36_249 ();
 fill_1 FILLER_36_251 ();
 decap_12 FILLER_36_253 ();
 decap_12 FILLER_36_265 ();
 decap_12 FILLER_36_277 ();
 decap_12 FILLER_36_289 ();
 fill_4 FILLER_36_301 ();
 fill_2 FILLER_36_305 ();
 fill_1 FILLER_36_307 ();
 decap_12 FILLER_36_309 ();
 decap_12 FILLER_36_321 ();
 decap_12 FILLER_36_333 ();
 decap_12 FILLER_36_345 ();
 fill_4 FILLER_36_357 ();
 fill_2 FILLER_36_361 ();
 fill_1 FILLER_36_363 ();
 decap_12 FILLER_36_365 ();
 decap_12 FILLER_36_377 ();
 decap_12 FILLER_36_389 ();
 decap_12 FILLER_36_401 ();
 fill_4 FILLER_36_413 ();
 fill_2 FILLER_36_417 ();
 fill_1 FILLER_36_419 ();
 decap_12 FILLER_36_421 ();
 decap_12 FILLER_36_433 ();
 decap_12 FILLER_36_445 ();
 decap_12 FILLER_36_457 ();
 fill_4 FILLER_36_469 ();
 fill_2 FILLER_36_473 ();
 fill_1 FILLER_36_475 ();
 decap_12 FILLER_36_477 ();
 decap_12 FILLER_36_489 ();
 decap_12 FILLER_36_501 ();
 decap_12 FILLER_36_513 ();
 fill_4 FILLER_36_525 ();
 fill_2 FILLER_36_529 ();
 fill_1 FILLER_36_531 ();
 decap_12 FILLER_36_533 ();
 decap_12 FILLER_36_545 ();
 decap_12 FILLER_36_557 ();
 decap_12 FILLER_36_569 ();
 fill_4 FILLER_36_581 ();
 fill_2 FILLER_36_585 ();
 fill_1 FILLER_36_587 ();
 decap_12 FILLER_36_589 ();
 decap_12 FILLER_36_601 ();
 decap_12 FILLER_36_613 ();
 decap_12 FILLER_37_3 ();
 decap_12 FILLER_37_15 ();
 decap_12 FILLER_37_27 ();
 decap_12 FILLER_37_39 ();
 fill_4 FILLER_37_51 ();
 fill_1 FILLER_37_55 ();
 decap_12 FILLER_37_57 ();
 decap_12 FILLER_37_69 ();
 decap_12 FILLER_37_81 ();
 decap_12 FILLER_37_93 ();
 fill_4 FILLER_37_105 ();
 fill_2 FILLER_37_109 ();
 fill_1 FILLER_37_111 ();
 decap_12 FILLER_37_113 ();
 decap_12 FILLER_37_125 ();
 decap_12 FILLER_37_137 ();
 decap_12 FILLER_37_149 ();
 fill_4 FILLER_37_161 ();
 fill_2 FILLER_37_165 ();
 fill_1 FILLER_37_167 ();
 decap_12 FILLER_37_169 ();
 decap_12 FILLER_37_181 ();
 decap_12 FILLER_37_193 ();
 decap_12 FILLER_37_205 ();
 fill_4 FILLER_37_217 ();
 fill_2 FILLER_37_221 ();
 fill_1 FILLER_37_223 ();
 decap_12 FILLER_37_225 ();
 decap_12 FILLER_37_237 ();
 decap_12 FILLER_37_249 ();
 decap_12 FILLER_37_261 ();
 fill_4 FILLER_37_273 ();
 fill_2 FILLER_37_277 ();
 fill_1 FILLER_37_279 ();
 decap_12 FILLER_37_281 ();
 decap_12 FILLER_37_293 ();
 decap_12 FILLER_37_305 ();
 decap_12 FILLER_37_317 ();
 fill_4 FILLER_37_329 ();
 fill_2 FILLER_37_333 ();
 fill_1 FILLER_37_335 ();
 decap_12 FILLER_37_337 ();
 decap_12 FILLER_37_349 ();
 decap_12 FILLER_37_361 ();
 decap_12 FILLER_37_373 ();
 fill_4 FILLER_37_385 ();
 fill_2 FILLER_37_389 ();
 fill_1 FILLER_37_391 ();
 decap_12 FILLER_37_393 ();
 decap_12 FILLER_37_405 ();
 decap_12 FILLER_37_417 ();
 decap_12 FILLER_37_429 ();
 fill_4 FILLER_37_441 ();
 fill_2 FILLER_37_445 ();
 fill_1 FILLER_37_447 ();
 decap_12 FILLER_37_449 ();
 decap_12 FILLER_37_461 ();
 decap_12 FILLER_37_473 ();
 decap_12 FILLER_37_485 ();
 fill_4 FILLER_37_497 ();
 fill_2 FILLER_37_501 ();
 fill_1 FILLER_37_503 ();
 decap_12 FILLER_37_505 ();
 decap_12 FILLER_37_517 ();
 decap_12 FILLER_37_529 ();
 decap_12 FILLER_37_541 ();
 fill_4 FILLER_37_553 ();
 fill_2 FILLER_37_557 ();
 fill_1 FILLER_37_559 ();
 decap_12 FILLER_37_561 ();
 decap_12 FILLER_37_573 ();
 decap_12 FILLER_37_585 ();
 decap_12 FILLER_37_597 ();
 fill_4 FILLER_37_609 ();
 fill_2 FILLER_37_613 ();
 fill_1 FILLER_37_615 ();
 fill_8 FILLER_37_617 ();
 decap_12 FILLER_38_3 ();
 decap_12 FILLER_38_15 ();
 fill_1 FILLER_38_27 ();
 decap_12 FILLER_38_29 ();
 decap_12 FILLER_38_41 ();
 decap_12 FILLER_38_53 ();
 decap_12 FILLER_38_65 ();
 fill_4 FILLER_38_77 ();
 fill_2 FILLER_38_81 ();
 fill_1 FILLER_38_83 ();
 decap_12 FILLER_38_85 ();
 decap_12 FILLER_38_97 ();
 decap_12 FILLER_38_109 ();
 decap_12 FILLER_38_121 ();
 fill_4 FILLER_38_133 ();
 fill_2 FILLER_38_137 ();
 fill_1 FILLER_38_139 ();
 decap_12 FILLER_38_141 ();
 decap_12 FILLER_38_153 ();
 decap_12 FILLER_38_165 ();
 decap_12 FILLER_38_177 ();
 fill_4 FILLER_38_189 ();
 fill_2 FILLER_38_193 ();
 fill_1 FILLER_38_195 ();
 decap_12 FILLER_38_197 ();
 decap_12 FILLER_38_209 ();
 decap_12 FILLER_38_221 ();
 decap_12 FILLER_38_233 ();
 fill_4 FILLER_38_245 ();
 fill_2 FILLER_38_249 ();
 fill_1 FILLER_38_251 ();
 decap_12 FILLER_38_253 ();
 decap_12 FILLER_38_265 ();
 decap_12 FILLER_38_277 ();
 decap_12 FILLER_38_289 ();
 fill_4 FILLER_38_301 ();
 fill_2 FILLER_38_305 ();
 fill_1 FILLER_38_307 ();
 decap_12 FILLER_38_309 ();
 decap_12 FILLER_38_321 ();
 decap_12 FILLER_38_333 ();
 decap_12 FILLER_38_345 ();
 fill_4 FILLER_38_357 ();
 fill_2 FILLER_38_361 ();
 fill_1 FILLER_38_363 ();
 decap_12 FILLER_38_365 ();
 decap_12 FILLER_38_377 ();
 decap_12 FILLER_38_389 ();
 decap_12 FILLER_38_401 ();
 fill_4 FILLER_38_413 ();
 fill_2 FILLER_38_417 ();
 fill_1 FILLER_38_419 ();
 decap_12 FILLER_38_421 ();
 decap_12 FILLER_38_433 ();
 decap_12 FILLER_38_445 ();
 decap_12 FILLER_38_457 ();
 fill_4 FILLER_38_469 ();
 fill_2 FILLER_38_473 ();
 fill_1 FILLER_38_475 ();
 decap_12 FILLER_38_477 ();
 decap_12 FILLER_38_489 ();
 decap_12 FILLER_38_501 ();
 decap_12 FILLER_38_513 ();
 fill_4 FILLER_38_525 ();
 fill_2 FILLER_38_529 ();
 fill_1 FILLER_38_531 ();
 decap_12 FILLER_38_533 ();
 decap_12 FILLER_38_545 ();
 decap_12 FILLER_38_557 ();
 decap_12 FILLER_38_569 ();
 fill_4 FILLER_38_581 ();
 fill_2 FILLER_38_585 ();
 fill_1 FILLER_38_587 ();
 decap_12 FILLER_38_589 ();
 decap_12 FILLER_38_601 ();
 decap_12 FILLER_38_613 ();
 decap_12 FILLER_39_3 ();
 decap_12 FILLER_39_15 ();
 decap_12 FILLER_39_27 ();
 decap_12 FILLER_39_39 ();
 fill_4 FILLER_39_51 ();
 fill_1 FILLER_39_55 ();
 decap_12 FILLER_39_57 ();
 decap_12 FILLER_39_69 ();
 decap_12 FILLER_39_81 ();
 decap_12 FILLER_39_93 ();
 fill_4 FILLER_39_105 ();
 fill_2 FILLER_39_109 ();
 fill_1 FILLER_39_111 ();
 decap_12 FILLER_39_113 ();
 decap_12 FILLER_39_125 ();
 decap_12 FILLER_39_137 ();
 decap_12 FILLER_39_149 ();
 fill_4 FILLER_39_161 ();
 fill_2 FILLER_39_165 ();
 fill_1 FILLER_39_167 ();
 decap_12 FILLER_39_169 ();
 decap_12 FILLER_39_181 ();
 decap_12 FILLER_39_193 ();
 decap_12 FILLER_39_205 ();
 fill_4 FILLER_39_217 ();
 fill_2 FILLER_39_221 ();
 fill_1 FILLER_39_223 ();
 decap_12 FILLER_39_225 ();
 decap_12 FILLER_39_237 ();
 decap_12 FILLER_39_249 ();
 decap_12 FILLER_39_261 ();
 fill_4 FILLER_39_273 ();
 fill_2 FILLER_39_277 ();
 fill_1 FILLER_39_279 ();
 decap_12 FILLER_39_281 ();
 decap_12 FILLER_39_293 ();
 decap_12 FILLER_39_305 ();
 decap_12 FILLER_39_317 ();
 fill_4 FILLER_39_329 ();
 fill_2 FILLER_39_333 ();
 fill_1 FILLER_39_335 ();
 decap_12 FILLER_39_337 ();
 decap_12 FILLER_39_349 ();
 decap_12 FILLER_39_361 ();
 decap_12 FILLER_39_373 ();
 fill_4 FILLER_39_385 ();
 fill_2 FILLER_39_389 ();
 fill_1 FILLER_39_391 ();
 decap_12 FILLER_39_393 ();
 decap_12 FILLER_39_405 ();
 decap_12 FILLER_39_417 ();
 decap_12 FILLER_39_429 ();
 fill_4 FILLER_39_441 ();
 fill_2 FILLER_39_445 ();
 fill_1 FILLER_39_447 ();
 decap_12 FILLER_39_449 ();
 decap_12 FILLER_39_461 ();
 decap_12 FILLER_39_473 ();
 decap_12 FILLER_39_485 ();
 fill_4 FILLER_39_497 ();
 fill_2 FILLER_39_501 ();
 fill_1 FILLER_39_503 ();
 decap_12 FILLER_39_505 ();
 decap_12 FILLER_39_517 ();
 decap_12 FILLER_39_529 ();
 decap_12 FILLER_39_541 ();
 fill_4 FILLER_39_553 ();
 fill_2 FILLER_39_557 ();
 fill_1 FILLER_39_559 ();
 decap_12 FILLER_39_561 ();
 decap_12 FILLER_39_573 ();
 decap_12 FILLER_39_585 ();
 decap_12 FILLER_39_597 ();
 fill_4 FILLER_39_609 ();
 fill_2 FILLER_39_613 ();
 fill_1 FILLER_39_615 ();
 fill_8 FILLER_39_617 ();
 decap_12 FILLER_40_3 ();
 decap_12 FILLER_40_15 ();
 fill_1 FILLER_40_27 ();
 decap_12 FILLER_40_29 ();
 decap_12 FILLER_40_41 ();
 decap_12 FILLER_40_53 ();
 decap_12 FILLER_40_65 ();
 fill_4 FILLER_40_77 ();
 fill_2 FILLER_40_81 ();
 fill_1 FILLER_40_83 ();
 decap_12 FILLER_40_85 ();
 decap_12 FILLER_40_97 ();
 decap_12 FILLER_40_109 ();
 decap_12 FILLER_40_121 ();
 fill_4 FILLER_40_133 ();
 fill_2 FILLER_40_137 ();
 fill_1 FILLER_40_139 ();
 decap_12 FILLER_40_141 ();
 decap_12 FILLER_40_153 ();
 decap_12 FILLER_40_165 ();
 decap_12 FILLER_40_177 ();
 fill_4 FILLER_40_189 ();
 fill_2 FILLER_40_193 ();
 fill_1 FILLER_40_195 ();
 decap_12 FILLER_40_197 ();
 decap_12 FILLER_40_209 ();
 decap_12 FILLER_40_221 ();
 decap_12 FILLER_40_233 ();
 fill_4 FILLER_40_245 ();
 fill_2 FILLER_40_249 ();
 fill_1 FILLER_40_251 ();
 decap_12 FILLER_40_253 ();
 decap_12 FILLER_40_265 ();
 decap_12 FILLER_40_277 ();
 decap_12 FILLER_40_289 ();
 fill_4 FILLER_40_301 ();
 fill_2 FILLER_40_305 ();
 fill_1 FILLER_40_307 ();
 decap_12 FILLER_40_309 ();
 decap_12 FILLER_40_321 ();
 decap_12 FILLER_40_333 ();
 decap_12 FILLER_40_345 ();
 fill_4 FILLER_40_357 ();
 fill_2 FILLER_40_361 ();
 fill_1 FILLER_40_363 ();
 decap_12 FILLER_40_365 ();
 decap_12 FILLER_40_377 ();
 decap_12 FILLER_40_389 ();
 decap_12 FILLER_40_401 ();
 fill_4 FILLER_40_413 ();
 fill_2 FILLER_40_417 ();
 fill_1 FILLER_40_419 ();
 decap_12 FILLER_40_421 ();
 decap_12 FILLER_40_433 ();
 decap_12 FILLER_40_445 ();
 decap_12 FILLER_40_457 ();
 fill_4 FILLER_40_469 ();
 fill_2 FILLER_40_473 ();
 fill_1 FILLER_40_475 ();
 decap_12 FILLER_40_477 ();
 decap_12 FILLER_40_489 ();
 decap_12 FILLER_40_501 ();
 decap_12 FILLER_40_513 ();
 fill_4 FILLER_40_525 ();
 fill_2 FILLER_40_529 ();
 fill_1 FILLER_40_531 ();
 decap_12 FILLER_40_533 ();
 decap_12 FILLER_40_545 ();
 decap_12 FILLER_40_557 ();
 decap_12 FILLER_40_569 ();
 fill_4 FILLER_40_581 ();
 fill_2 FILLER_40_585 ();
 fill_1 FILLER_40_587 ();
 decap_12 FILLER_40_589 ();
 decap_12 FILLER_40_601 ();
 decap_12 FILLER_40_613 ();
 decap_12 FILLER_41_3 ();
 decap_12 FILLER_41_15 ();
 decap_12 FILLER_41_27 ();
 decap_12 FILLER_41_39 ();
 fill_4 FILLER_41_51 ();
 fill_1 FILLER_41_55 ();
 decap_12 FILLER_41_57 ();
 decap_12 FILLER_41_69 ();
 decap_12 FILLER_41_81 ();
 decap_12 FILLER_41_93 ();
 fill_4 FILLER_41_105 ();
 fill_2 FILLER_41_109 ();
 fill_1 FILLER_41_111 ();
 decap_12 FILLER_41_113 ();
 decap_12 FILLER_41_125 ();
 decap_12 FILLER_41_137 ();
 decap_12 FILLER_41_149 ();
 fill_4 FILLER_41_161 ();
 fill_2 FILLER_41_165 ();
 fill_1 FILLER_41_167 ();
 decap_12 FILLER_41_169 ();
 decap_12 FILLER_41_181 ();
 decap_12 FILLER_41_193 ();
 decap_12 FILLER_41_205 ();
 fill_4 FILLER_41_217 ();
 fill_2 FILLER_41_221 ();
 fill_1 FILLER_41_223 ();
 decap_12 FILLER_41_225 ();
 decap_12 FILLER_41_237 ();
 decap_12 FILLER_41_249 ();
 decap_12 FILLER_41_261 ();
 fill_4 FILLER_41_273 ();
 fill_2 FILLER_41_277 ();
 fill_1 FILLER_41_279 ();
 decap_12 FILLER_41_281 ();
 decap_12 FILLER_41_293 ();
 decap_12 FILLER_41_305 ();
 decap_12 FILLER_41_317 ();
 fill_4 FILLER_41_329 ();
 fill_2 FILLER_41_333 ();
 fill_1 FILLER_41_335 ();
 decap_12 FILLER_41_337 ();
 decap_12 FILLER_41_349 ();
 decap_12 FILLER_41_361 ();
 decap_12 FILLER_41_373 ();
 fill_4 FILLER_41_385 ();
 fill_2 FILLER_41_389 ();
 fill_1 FILLER_41_391 ();
 decap_12 FILLER_41_393 ();
 decap_12 FILLER_41_405 ();
 decap_12 FILLER_41_417 ();
 decap_12 FILLER_41_429 ();
 fill_4 FILLER_41_441 ();
 fill_2 FILLER_41_445 ();
 fill_1 FILLER_41_447 ();
 decap_12 FILLER_41_449 ();
 decap_12 FILLER_41_461 ();
 decap_12 FILLER_41_473 ();
 decap_12 FILLER_41_485 ();
 fill_4 FILLER_41_497 ();
 fill_2 FILLER_41_501 ();
 fill_1 FILLER_41_503 ();
 decap_12 FILLER_41_505 ();
 decap_12 FILLER_41_517 ();
 decap_12 FILLER_41_529 ();
 decap_12 FILLER_41_541 ();
 fill_4 FILLER_41_553 ();
 fill_2 FILLER_41_557 ();
 fill_1 FILLER_41_559 ();
 decap_12 FILLER_41_561 ();
 decap_12 FILLER_41_573 ();
 decap_12 FILLER_41_585 ();
 decap_12 FILLER_41_597 ();
 fill_4 FILLER_41_609 ();
 fill_2 FILLER_41_613 ();
 fill_1 FILLER_41_615 ();
 fill_8 FILLER_41_617 ();
 decap_12 FILLER_42_3 ();
 decap_12 FILLER_42_15 ();
 fill_1 FILLER_42_27 ();
 decap_12 FILLER_42_29 ();
 decap_12 FILLER_42_41 ();
 decap_12 FILLER_42_53 ();
 decap_12 FILLER_42_65 ();
 fill_4 FILLER_42_77 ();
 fill_2 FILLER_42_81 ();
 fill_1 FILLER_42_83 ();
 decap_12 FILLER_42_85 ();
 decap_12 FILLER_42_97 ();
 decap_12 FILLER_42_109 ();
 decap_12 FILLER_42_121 ();
 fill_4 FILLER_42_133 ();
 fill_2 FILLER_42_137 ();
 fill_1 FILLER_42_139 ();
 decap_12 FILLER_42_141 ();
 decap_12 FILLER_42_153 ();
 decap_12 FILLER_42_165 ();
 decap_12 FILLER_42_177 ();
 fill_4 FILLER_42_189 ();
 fill_2 FILLER_42_193 ();
 fill_1 FILLER_42_195 ();
 decap_12 FILLER_42_197 ();
 decap_12 FILLER_42_209 ();
 decap_12 FILLER_42_221 ();
 decap_12 FILLER_42_233 ();
 fill_4 FILLER_42_245 ();
 fill_2 FILLER_42_249 ();
 fill_1 FILLER_42_251 ();
 decap_12 FILLER_42_253 ();
 decap_12 FILLER_42_265 ();
 decap_12 FILLER_42_277 ();
 decap_12 FILLER_42_289 ();
 fill_4 FILLER_42_301 ();
 fill_2 FILLER_42_305 ();
 fill_1 FILLER_42_307 ();
 decap_12 FILLER_42_309 ();
 decap_12 FILLER_42_321 ();
 decap_12 FILLER_42_333 ();
 decap_12 FILLER_42_345 ();
 fill_4 FILLER_42_357 ();
 fill_2 FILLER_42_361 ();
 fill_1 FILLER_42_363 ();
 decap_12 FILLER_42_365 ();
 decap_12 FILLER_42_377 ();
 decap_12 FILLER_42_389 ();
 decap_12 FILLER_42_401 ();
 fill_4 FILLER_42_413 ();
 fill_2 FILLER_42_417 ();
 fill_1 FILLER_42_419 ();
 decap_12 FILLER_42_421 ();
 decap_12 FILLER_42_433 ();
 decap_12 FILLER_42_445 ();
 decap_12 FILLER_42_457 ();
 fill_4 FILLER_42_469 ();
 fill_2 FILLER_42_473 ();
 fill_1 FILLER_42_475 ();
 decap_12 FILLER_42_477 ();
 decap_12 FILLER_42_489 ();
 decap_12 FILLER_42_501 ();
 decap_12 FILLER_42_513 ();
 fill_4 FILLER_42_525 ();
 fill_2 FILLER_42_529 ();
 fill_1 FILLER_42_531 ();
 decap_12 FILLER_42_533 ();
 decap_12 FILLER_42_545 ();
 decap_12 FILLER_42_557 ();
 decap_12 FILLER_42_569 ();
 fill_4 FILLER_42_581 ();
 fill_2 FILLER_42_585 ();
 fill_1 FILLER_42_587 ();
 decap_12 FILLER_42_589 ();
 decap_12 FILLER_42_601 ();
 decap_12 FILLER_42_613 ();
 decap_12 FILLER_43_3 ();
 decap_12 FILLER_43_15 ();
 decap_12 FILLER_43_27 ();
 decap_12 FILLER_43_39 ();
 fill_4 FILLER_43_51 ();
 fill_1 FILLER_43_55 ();
 decap_12 FILLER_43_57 ();
 decap_12 FILLER_43_69 ();
 decap_12 FILLER_43_81 ();
 decap_12 FILLER_43_93 ();
 fill_4 FILLER_43_105 ();
 fill_2 FILLER_43_109 ();
 fill_1 FILLER_43_111 ();
 decap_12 FILLER_43_113 ();
 decap_12 FILLER_43_125 ();
 decap_12 FILLER_43_137 ();
 decap_12 FILLER_43_149 ();
 fill_4 FILLER_43_161 ();
 fill_2 FILLER_43_165 ();
 fill_1 FILLER_43_167 ();
 decap_12 FILLER_43_169 ();
 decap_12 FILLER_43_181 ();
 decap_12 FILLER_43_193 ();
 decap_12 FILLER_43_205 ();
 fill_4 FILLER_43_217 ();
 fill_2 FILLER_43_221 ();
 fill_1 FILLER_43_223 ();
 decap_12 FILLER_43_225 ();
 decap_12 FILLER_43_237 ();
 decap_12 FILLER_43_249 ();
 decap_12 FILLER_43_261 ();
 fill_4 FILLER_43_273 ();
 fill_2 FILLER_43_277 ();
 fill_1 FILLER_43_279 ();
 decap_12 FILLER_43_281 ();
 decap_12 FILLER_43_293 ();
 decap_12 FILLER_43_305 ();
 decap_12 FILLER_43_317 ();
 fill_4 FILLER_43_329 ();
 fill_2 FILLER_43_333 ();
 fill_1 FILLER_43_335 ();
 decap_12 FILLER_43_337 ();
 decap_12 FILLER_43_349 ();
 decap_12 FILLER_43_361 ();
 decap_12 FILLER_43_373 ();
 fill_4 FILLER_43_385 ();
 fill_2 FILLER_43_389 ();
 fill_1 FILLER_43_391 ();
 decap_12 FILLER_43_393 ();
 decap_12 FILLER_43_405 ();
 decap_12 FILLER_43_417 ();
 decap_12 FILLER_43_429 ();
 fill_4 FILLER_43_441 ();
 fill_2 FILLER_43_445 ();
 fill_1 FILLER_43_447 ();
 decap_12 FILLER_43_449 ();
 decap_12 FILLER_43_461 ();
 decap_12 FILLER_43_473 ();
 decap_12 FILLER_43_485 ();
 fill_4 FILLER_43_497 ();
 fill_2 FILLER_43_501 ();
 fill_1 FILLER_43_503 ();
 decap_12 FILLER_43_505 ();
 decap_12 FILLER_43_517 ();
 decap_12 FILLER_43_529 ();
 decap_12 FILLER_43_541 ();
 fill_4 FILLER_43_553 ();
 fill_2 FILLER_43_557 ();
 fill_1 FILLER_43_559 ();
 decap_12 FILLER_43_561 ();
 decap_12 FILLER_43_573 ();
 decap_12 FILLER_43_585 ();
 decap_12 FILLER_43_597 ();
 fill_4 FILLER_43_609 ();
 fill_2 FILLER_43_613 ();
 fill_1 FILLER_43_615 ();
 fill_8 FILLER_43_617 ();
 decap_12 FILLER_44_3 ();
 decap_12 FILLER_44_15 ();
 fill_1 FILLER_44_27 ();
 decap_12 FILLER_44_29 ();
 decap_12 FILLER_44_41 ();
 decap_12 FILLER_44_53 ();
 decap_12 FILLER_44_65 ();
 fill_4 FILLER_44_77 ();
 fill_2 FILLER_44_81 ();
 fill_1 FILLER_44_83 ();
 decap_12 FILLER_44_85 ();
 decap_12 FILLER_44_97 ();
 decap_12 FILLER_44_109 ();
 decap_12 FILLER_44_121 ();
 fill_4 FILLER_44_133 ();
 fill_2 FILLER_44_137 ();
 fill_1 FILLER_44_139 ();
 decap_12 FILLER_44_141 ();
 decap_12 FILLER_44_153 ();
 decap_12 FILLER_44_165 ();
 decap_12 FILLER_44_177 ();
 fill_4 FILLER_44_189 ();
 fill_2 FILLER_44_193 ();
 fill_1 FILLER_44_195 ();
 decap_12 FILLER_44_197 ();
 decap_12 FILLER_44_209 ();
 decap_12 FILLER_44_221 ();
 decap_12 FILLER_44_233 ();
 fill_4 FILLER_44_245 ();
 fill_2 FILLER_44_249 ();
 fill_1 FILLER_44_251 ();
 decap_12 FILLER_44_253 ();
 decap_12 FILLER_44_265 ();
 decap_12 FILLER_44_277 ();
 decap_12 FILLER_44_289 ();
 fill_4 FILLER_44_301 ();
 fill_2 FILLER_44_305 ();
 fill_1 FILLER_44_307 ();
 decap_12 FILLER_44_309 ();
 decap_12 FILLER_44_321 ();
 decap_12 FILLER_44_333 ();
 decap_12 FILLER_44_345 ();
 fill_4 FILLER_44_357 ();
 fill_2 FILLER_44_361 ();
 fill_1 FILLER_44_363 ();
 decap_12 FILLER_44_365 ();
 decap_12 FILLER_44_377 ();
 decap_12 FILLER_44_389 ();
 decap_12 FILLER_44_401 ();
 fill_4 FILLER_44_413 ();
 fill_2 FILLER_44_417 ();
 fill_1 FILLER_44_419 ();
 decap_12 FILLER_44_421 ();
 decap_12 FILLER_44_433 ();
 decap_12 FILLER_44_445 ();
 decap_12 FILLER_44_457 ();
 fill_4 FILLER_44_469 ();
 fill_2 FILLER_44_473 ();
 fill_1 FILLER_44_475 ();
 decap_12 FILLER_44_477 ();
 decap_12 FILLER_44_489 ();
 decap_12 FILLER_44_501 ();
 decap_12 FILLER_44_513 ();
 fill_4 FILLER_44_525 ();
 fill_2 FILLER_44_529 ();
 fill_1 FILLER_44_531 ();
 decap_12 FILLER_44_533 ();
 decap_12 FILLER_44_545 ();
 decap_12 FILLER_44_557 ();
 decap_12 FILLER_44_569 ();
 fill_4 FILLER_44_581 ();
 fill_2 FILLER_44_585 ();
 fill_1 FILLER_44_587 ();
 decap_12 FILLER_44_589 ();
 decap_12 FILLER_44_601 ();
 decap_12 FILLER_44_613 ();
 decap_12 FILLER_45_3 ();
 decap_12 FILLER_45_15 ();
 decap_12 FILLER_45_27 ();
 decap_12 FILLER_45_39 ();
 fill_4 FILLER_45_51 ();
 fill_1 FILLER_45_55 ();
 decap_12 FILLER_45_57 ();
 decap_12 FILLER_45_69 ();
 decap_12 FILLER_45_81 ();
 decap_12 FILLER_45_93 ();
 fill_4 FILLER_45_105 ();
 fill_2 FILLER_45_109 ();
 fill_1 FILLER_45_111 ();
 decap_12 FILLER_45_113 ();
 decap_12 FILLER_45_125 ();
 decap_12 FILLER_45_137 ();
 decap_12 FILLER_45_149 ();
 fill_4 FILLER_45_161 ();
 fill_2 FILLER_45_165 ();
 fill_1 FILLER_45_167 ();
 decap_12 FILLER_45_169 ();
 decap_12 FILLER_45_181 ();
 decap_12 FILLER_45_193 ();
 decap_12 FILLER_45_205 ();
 fill_4 FILLER_45_217 ();
 fill_2 FILLER_45_221 ();
 fill_1 FILLER_45_223 ();
 decap_12 FILLER_45_225 ();
 decap_12 FILLER_45_237 ();
 decap_12 FILLER_45_249 ();
 decap_12 FILLER_45_261 ();
 fill_4 FILLER_45_273 ();
 fill_2 FILLER_45_277 ();
 fill_1 FILLER_45_279 ();
 decap_12 FILLER_45_281 ();
 decap_12 FILLER_45_293 ();
 decap_12 FILLER_45_305 ();
 decap_12 FILLER_45_317 ();
 fill_4 FILLER_45_329 ();
 fill_2 FILLER_45_333 ();
 fill_1 FILLER_45_335 ();
 decap_12 FILLER_45_337 ();
 decap_12 FILLER_45_349 ();
 decap_12 FILLER_45_361 ();
 decap_12 FILLER_45_373 ();
 fill_4 FILLER_45_385 ();
 fill_2 FILLER_45_389 ();
 fill_1 FILLER_45_391 ();
 decap_12 FILLER_45_393 ();
 decap_12 FILLER_45_405 ();
 decap_12 FILLER_45_417 ();
 decap_12 FILLER_45_429 ();
 fill_4 FILLER_45_441 ();
 fill_2 FILLER_45_445 ();
 fill_1 FILLER_45_447 ();
 decap_12 FILLER_45_449 ();
 decap_12 FILLER_45_461 ();
 decap_12 FILLER_45_473 ();
 decap_12 FILLER_45_485 ();
 fill_4 FILLER_45_497 ();
 fill_2 FILLER_45_501 ();
 fill_1 FILLER_45_503 ();
 decap_12 FILLER_45_505 ();
 decap_12 FILLER_45_517 ();
 decap_12 FILLER_45_529 ();
 decap_12 FILLER_45_541 ();
 fill_4 FILLER_45_553 ();
 fill_2 FILLER_45_557 ();
 fill_1 FILLER_45_559 ();
 decap_12 FILLER_45_561 ();
 decap_12 FILLER_45_573 ();
 decap_12 FILLER_45_585 ();
 decap_12 FILLER_45_597 ();
 fill_4 FILLER_45_609 ();
 fill_2 FILLER_45_613 ();
 fill_1 FILLER_45_615 ();
 fill_8 FILLER_45_617 ();
 decap_12 FILLER_46_3 ();
 decap_12 FILLER_46_15 ();
 fill_1 FILLER_46_27 ();
 decap_12 FILLER_46_29 ();
 decap_12 FILLER_46_41 ();
 decap_12 FILLER_46_53 ();
 decap_12 FILLER_46_65 ();
 fill_4 FILLER_46_77 ();
 fill_2 FILLER_46_81 ();
 fill_1 FILLER_46_83 ();
 decap_12 FILLER_46_85 ();
 decap_12 FILLER_46_97 ();
 decap_12 FILLER_46_109 ();
 decap_12 FILLER_46_121 ();
 fill_4 FILLER_46_133 ();
 fill_2 FILLER_46_137 ();
 fill_1 FILLER_46_139 ();
 decap_12 FILLER_46_141 ();
 decap_12 FILLER_46_153 ();
 decap_12 FILLER_46_165 ();
 decap_12 FILLER_46_177 ();
 fill_4 FILLER_46_189 ();
 fill_2 FILLER_46_193 ();
 fill_1 FILLER_46_195 ();
 decap_12 FILLER_46_197 ();
 decap_12 FILLER_46_209 ();
 decap_12 FILLER_46_221 ();
 decap_12 FILLER_46_233 ();
 fill_4 FILLER_46_245 ();
 fill_2 FILLER_46_249 ();
 fill_1 FILLER_46_251 ();
 decap_12 FILLER_46_253 ();
 decap_12 FILLER_46_265 ();
 decap_12 FILLER_46_277 ();
 decap_12 FILLER_46_289 ();
 fill_4 FILLER_46_301 ();
 fill_2 FILLER_46_305 ();
 fill_1 FILLER_46_307 ();
 decap_12 FILLER_46_309 ();
 decap_12 FILLER_46_321 ();
 decap_12 FILLER_46_333 ();
 decap_12 FILLER_46_345 ();
 fill_4 FILLER_46_357 ();
 fill_2 FILLER_46_361 ();
 fill_1 FILLER_46_363 ();
 decap_12 FILLER_46_365 ();
 decap_12 FILLER_46_377 ();
 decap_12 FILLER_46_389 ();
 decap_12 FILLER_46_401 ();
 fill_4 FILLER_46_413 ();
 fill_2 FILLER_46_417 ();
 fill_1 FILLER_46_419 ();
 decap_12 FILLER_46_421 ();
 decap_12 FILLER_46_433 ();
 decap_12 FILLER_46_445 ();
 decap_12 FILLER_46_457 ();
 fill_4 FILLER_46_469 ();
 fill_2 FILLER_46_473 ();
 fill_1 FILLER_46_475 ();
 decap_12 FILLER_46_477 ();
 decap_12 FILLER_46_489 ();
 decap_12 FILLER_46_501 ();
 decap_12 FILLER_46_513 ();
 fill_4 FILLER_46_525 ();
 fill_2 FILLER_46_529 ();
 fill_1 FILLER_46_531 ();
 decap_12 FILLER_46_533 ();
 decap_12 FILLER_46_545 ();
 decap_12 FILLER_46_557 ();
 decap_12 FILLER_46_569 ();
 fill_4 FILLER_46_581 ();
 fill_2 FILLER_46_585 ();
 fill_1 FILLER_46_587 ();
 decap_12 FILLER_46_589 ();
 decap_12 FILLER_46_601 ();
 decap_12 FILLER_46_613 ();
 decap_12 FILLER_47_3 ();
 decap_12 FILLER_47_15 ();
 decap_12 FILLER_47_27 ();
 decap_12 FILLER_47_39 ();
 fill_4 FILLER_47_51 ();
 fill_1 FILLER_47_55 ();
 decap_12 FILLER_47_57 ();
 decap_12 FILLER_47_69 ();
 decap_12 FILLER_47_81 ();
 decap_12 FILLER_47_93 ();
 fill_4 FILLER_47_105 ();
 fill_2 FILLER_47_109 ();
 fill_1 FILLER_47_111 ();
 decap_12 FILLER_47_113 ();
 decap_12 FILLER_47_125 ();
 decap_12 FILLER_47_137 ();
 decap_12 FILLER_47_149 ();
 fill_4 FILLER_47_161 ();
 fill_2 FILLER_47_165 ();
 fill_1 FILLER_47_167 ();
 decap_12 FILLER_47_169 ();
 decap_12 FILLER_47_181 ();
 decap_12 FILLER_47_193 ();
 decap_12 FILLER_47_205 ();
 fill_4 FILLER_47_217 ();
 fill_2 FILLER_47_221 ();
 fill_1 FILLER_47_223 ();
 decap_12 FILLER_47_225 ();
 decap_12 FILLER_47_237 ();
 decap_12 FILLER_47_249 ();
 decap_12 FILLER_47_261 ();
 fill_4 FILLER_47_273 ();
 fill_2 FILLER_47_277 ();
 fill_1 FILLER_47_279 ();
 decap_12 FILLER_47_281 ();
 decap_12 FILLER_47_293 ();
 decap_12 FILLER_47_305 ();
 decap_12 FILLER_47_317 ();
 fill_4 FILLER_47_329 ();
 fill_2 FILLER_47_333 ();
 fill_1 FILLER_47_335 ();
 decap_12 FILLER_47_337 ();
 decap_12 FILLER_47_349 ();
 decap_12 FILLER_47_361 ();
 decap_12 FILLER_47_373 ();
 fill_4 FILLER_47_385 ();
 fill_2 FILLER_47_389 ();
 fill_1 FILLER_47_391 ();
 decap_12 FILLER_47_393 ();
 decap_12 FILLER_47_405 ();
 decap_12 FILLER_47_417 ();
 decap_12 FILLER_47_429 ();
 fill_4 FILLER_47_441 ();
 fill_2 FILLER_47_445 ();
 fill_1 FILLER_47_447 ();
 decap_12 FILLER_47_449 ();
 decap_12 FILLER_47_461 ();
 decap_12 FILLER_47_473 ();
 decap_12 FILLER_47_485 ();
 fill_4 FILLER_47_497 ();
 fill_2 FILLER_47_501 ();
 fill_1 FILLER_47_503 ();
 decap_12 FILLER_47_505 ();
 decap_12 FILLER_47_517 ();
 decap_12 FILLER_47_529 ();
 decap_12 FILLER_47_541 ();
 fill_4 FILLER_47_553 ();
 fill_2 FILLER_47_557 ();
 fill_1 FILLER_47_559 ();
 decap_12 FILLER_47_561 ();
 decap_12 FILLER_47_573 ();
 decap_12 FILLER_47_585 ();
 decap_12 FILLER_47_597 ();
 fill_4 FILLER_47_609 ();
 fill_2 FILLER_47_613 ();
 fill_1 FILLER_47_615 ();
 fill_8 FILLER_47_617 ();
 decap_12 FILLER_48_3 ();
 decap_12 FILLER_48_15 ();
 fill_1 FILLER_48_27 ();
 decap_12 FILLER_48_29 ();
 decap_12 FILLER_48_41 ();
 decap_12 FILLER_48_53 ();
 decap_12 FILLER_48_65 ();
 fill_4 FILLER_48_77 ();
 fill_2 FILLER_48_81 ();
 fill_1 FILLER_48_83 ();
 decap_12 FILLER_48_85 ();
 decap_12 FILLER_48_97 ();
 decap_12 FILLER_48_109 ();
 decap_12 FILLER_48_121 ();
 fill_4 FILLER_48_133 ();
 fill_2 FILLER_48_137 ();
 fill_1 FILLER_48_139 ();
 decap_12 FILLER_48_141 ();
 decap_12 FILLER_48_153 ();
 decap_12 FILLER_48_165 ();
 decap_12 FILLER_48_177 ();
 fill_4 FILLER_48_189 ();
 fill_2 FILLER_48_193 ();
 fill_1 FILLER_48_195 ();
 decap_12 FILLER_48_197 ();
 decap_12 FILLER_48_209 ();
 decap_12 FILLER_48_221 ();
 decap_12 FILLER_48_233 ();
 fill_4 FILLER_48_245 ();
 fill_2 FILLER_48_249 ();
 fill_1 FILLER_48_251 ();
 decap_12 FILLER_48_253 ();
 decap_12 FILLER_48_265 ();
 decap_12 FILLER_48_277 ();
 decap_12 FILLER_48_289 ();
 fill_4 FILLER_48_301 ();
 fill_2 FILLER_48_305 ();
 fill_1 FILLER_48_307 ();
 decap_12 FILLER_48_309 ();
 decap_12 FILLER_48_321 ();
 decap_12 FILLER_48_333 ();
 decap_12 FILLER_48_345 ();
 fill_4 FILLER_48_357 ();
 fill_2 FILLER_48_361 ();
 fill_1 FILLER_48_363 ();
 decap_12 FILLER_48_365 ();
 decap_12 FILLER_48_377 ();
 decap_12 FILLER_48_389 ();
 decap_12 FILLER_48_401 ();
 fill_4 FILLER_48_413 ();
 fill_2 FILLER_48_417 ();
 fill_1 FILLER_48_419 ();
 decap_12 FILLER_48_421 ();
 decap_12 FILLER_48_433 ();
 decap_12 FILLER_48_445 ();
 decap_12 FILLER_48_457 ();
 fill_4 FILLER_48_469 ();
 fill_2 FILLER_48_473 ();
 fill_1 FILLER_48_475 ();
 decap_12 FILLER_48_477 ();
 decap_12 FILLER_48_489 ();
 decap_12 FILLER_48_501 ();
 decap_12 FILLER_48_513 ();
 fill_4 FILLER_48_525 ();
 fill_2 FILLER_48_529 ();
 fill_1 FILLER_48_531 ();
 decap_12 FILLER_48_533 ();
 decap_12 FILLER_48_545 ();
 decap_12 FILLER_48_557 ();
 decap_12 FILLER_48_569 ();
 fill_4 FILLER_48_581 ();
 fill_2 FILLER_48_585 ();
 fill_1 FILLER_48_587 ();
 decap_12 FILLER_48_589 ();
 decap_12 FILLER_48_601 ();
 decap_12 FILLER_48_613 ();
 decap_12 FILLER_49_3 ();
 decap_12 FILLER_49_15 ();
 decap_12 FILLER_49_27 ();
 decap_12 FILLER_49_39 ();
 fill_4 FILLER_49_51 ();
 fill_1 FILLER_49_55 ();
 decap_12 FILLER_49_57 ();
 decap_12 FILLER_49_69 ();
 decap_12 FILLER_49_81 ();
 decap_12 FILLER_49_93 ();
 fill_4 FILLER_49_105 ();
 fill_2 FILLER_49_109 ();
 fill_1 FILLER_49_111 ();
 decap_12 FILLER_49_113 ();
 decap_12 FILLER_49_125 ();
 decap_12 FILLER_49_137 ();
 decap_12 FILLER_49_149 ();
 fill_4 FILLER_49_161 ();
 fill_2 FILLER_49_165 ();
 fill_1 FILLER_49_167 ();
 decap_12 FILLER_49_169 ();
 decap_12 FILLER_49_181 ();
 decap_12 FILLER_49_193 ();
 decap_12 FILLER_49_205 ();
 fill_4 FILLER_49_217 ();
 fill_2 FILLER_49_221 ();
 fill_1 FILLER_49_223 ();
 decap_12 FILLER_49_225 ();
 decap_12 FILLER_49_237 ();
 decap_12 FILLER_49_249 ();
 decap_12 FILLER_49_261 ();
 fill_4 FILLER_49_273 ();
 fill_2 FILLER_49_277 ();
 fill_1 FILLER_49_279 ();
 decap_12 FILLER_49_281 ();
 decap_12 FILLER_49_293 ();
 decap_12 FILLER_49_305 ();
 decap_12 FILLER_49_317 ();
 fill_4 FILLER_49_329 ();
 fill_2 FILLER_49_333 ();
 fill_1 FILLER_49_335 ();
 decap_12 FILLER_49_337 ();
 decap_12 FILLER_49_349 ();
 decap_12 FILLER_49_361 ();
 decap_12 FILLER_49_373 ();
 fill_4 FILLER_49_385 ();
 fill_2 FILLER_49_389 ();
 fill_1 FILLER_49_391 ();
 decap_12 FILLER_49_393 ();
 decap_12 FILLER_49_405 ();
 decap_12 FILLER_49_417 ();
 decap_12 FILLER_49_429 ();
 fill_4 FILLER_49_441 ();
 fill_2 FILLER_49_445 ();
 fill_1 FILLER_49_447 ();
 decap_12 FILLER_49_449 ();
 decap_12 FILLER_49_461 ();
 decap_12 FILLER_49_473 ();
 decap_12 FILLER_49_485 ();
 fill_4 FILLER_49_497 ();
 fill_2 FILLER_49_501 ();
 fill_1 FILLER_49_503 ();
 decap_12 FILLER_49_505 ();
 decap_12 FILLER_49_517 ();
 decap_12 FILLER_49_529 ();
 decap_12 FILLER_49_541 ();
 fill_4 FILLER_49_553 ();
 fill_2 FILLER_49_557 ();
 fill_1 FILLER_49_559 ();
 decap_12 FILLER_49_561 ();
 decap_12 FILLER_49_573 ();
 decap_12 FILLER_49_585 ();
 decap_12 FILLER_49_597 ();
 fill_4 FILLER_49_609 ();
 fill_2 FILLER_49_613 ();
 fill_1 FILLER_49_615 ();
 fill_8 FILLER_49_617 ();
 decap_12 FILLER_50_13 ();
 fill_2 FILLER_50_25 ();
 fill_1 FILLER_50_27 ();
 decap_12 FILLER_50_51 ();
 decap_12 FILLER_50_63 ();
 fill_8 FILLER_50_75 ();
 fill_1 FILLER_50_83 ();
 decap_12 FILLER_50_85 ();
 decap_12 FILLER_50_97 ();
 decap_12 FILLER_50_109 ();
 decap_12 FILLER_50_121 ();
 fill_4 FILLER_50_133 ();
 fill_2 FILLER_50_137 ();
 fill_1 FILLER_50_139 ();
 decap_12 FILLER_50_141 ();
 decap_12 FILLER_50_153 ();
 decap_12 FILLER_50_165 ();
 decap_12 FILLER_50_177 ();
 fill_4 FILLER_50_189 ();
 fill_2 FILLER_50_193 ();
 fill_1 FILLER_50_195 ();
 decap_12 FILLER_50_197 ();
 decap_12 FILLER_50_209 ();
 decap_12 FILLER_50_221 ();
 decap_12 FILLER_50_233 ();
 fill_4 FILLER_50_245 ();
 fill_2 FILLER_50_249 ();
 fill_1 FILLER_50_251 ();
 decap_12 FILLER_50_253 ();
 decap_12 FILLER_50_265 ();
 decap_12 FILLER_50_277 ();
 decap_12 FILLER_50_289 ();
 fill_4 FILLER_50_301 ();
 fill_2 FILLER_50_305 ();
 fill_1 FILLER_50_307 ();
 decap_12 FILLER_50_309 ();
 decap_12 FILLER_50_321 ();
 decap_12 FILLER_50_333 ();
 decap_12 FILLER_50_345 ();
 fill_4 FILLER_50_357 ();
 fill_2 FILLER_50_361 ();
 fill_1 FILLER_50_363 ();
 decap_12 FILLER_50_365 ();
 decap_12 FILLER_50_377 ();
 decap_12 FILLER_50_389 ();
 decap_12 FILLER_50_401 ();
 fill_4 FILLER_50_413 ();
 fill_2 FILLER_50_417 ();
 fill_1 FILLER_50_419 ();
 decap_12 FILLER_50_421 ();
 decap_12 FILLER_50_433 ();
 decap_12 FILLER_50_445 ();
 decap_12 FILLER_50_457 ();
 fill_4 FILLER_50_469 ();
 fill_2 FILLER_50_473 ();
 fill_1 FILLER_50_475 ();
 decap_12 FILLER_50_477 ();
 decap_12 FILLER_50_489 ();
 decap_12 FILLER_50_501 ();
 decap_12 FILLER_50_513 ();
 fill_4 FILLER_50_525 ();
 fill_2 FILLER_50_529 ();
 fill_1 FILLER_50_531 ();
 decap_12 FILLER_50_533 ();
 decap_12 FILLER_50_545 ();
 decap_12 FILLER_50_557 ();
 decap_12 FILLER_50_569 ();
 fill_4 FILLER_50_581 ();
 fill_2 FILLER_50_585 ();
 fill_1 FILLER_50_587 ();
 decap_12 FILLER_50_589 ();
 decap_12 FILLER_50_601 ();
 decap_12 FILLER_50_613 ();
 decap_12 FILLER_51_7 ();
 decap_12 FILLER_51_19 ();
 decap_12 FILLER_51_31 ();
 decap_12 FILLER_51_43 ();
 fill_1 FILLER_51_55 ();
 decap_12 FILLER_51_57 ();
 decap_12 FILLER_51_69 ();
 decap_12 FILLER_51_81 ();
 decap_12 FILLER_51_93 ();
 fill_4 FILLER_51_105 ();
 fill_2 FILLER_51_109 ();
 fill_1 FILLER_51_111 ();
 decap_12 FILLER_51_113 ();
 decap_12 FILLER_51_125 ();
 decap_12 FILLER_51_137 ();
 decap_12 FILLER_51_149 ();
 fill_4 FILLER_51_161 ();
 fill_2 FILLER_51_165 ();
 fill_1 FILLER_51_167 ();
 decap_12 FILLER_51_169 ();
 decap_12 FILLER_51_181 ();
 decap_12 FILLER_51_193 ();
 decap_12 FILLER_51_205 ();
 fill_4 FILLER_51_217 ();
 fill_2 FILLER_51_221 ();
 fill_1 FILLER_51_223 ();
 decap_12 FILLER_51_225 ();
 decap_12 FILLER_51_237 ();
 decap_12 FILLER_51_249 ();
 decap_12 FILLER_51_261 ();
 fill_4 FILLER_51_273 ();
 fill_2 FILLER_51_277 ();
 fill_1 FILLER_51_279 ();
 decap_12 FILLER_51_281 ();
 decap_12 FILLER_51_293 ();
 decap_12 FILLER_51_305 ();
 decap_12 FILLER_51_317 ();
 fill_4 FILLER_51_329 ();
 fill_2 FILLER_51_333 ();
 fill_1 FILLER_51_335 ();
 decap_12 FILLER_51_337 ();
 decap_12 FILLER_51_349 ();
 decap_12 FILLER_51_361 ();
 decap_12 FILLER_51_373 ();
 fill_4 FILLER_51_385 ();
 fill_2 FILLER_51_389 ();
 fill_1 FILLER_51_391 ();
 decap_12 FILLER_51_393 ();
 decap_12 FILLER_51_405 ();
 decap_12 FILLER_51_417 ();
 decap_12 FILLER_51_429 ();
 fill_4 FILLER_51_441 ();
 fill_2 FILLER_51_445 ();
 fill_1 FILLER_51_447 ();
 decap_12 FILLER_51_449 ();
 decap_12 FILLER_51_461 ();
 decap_12 FILLER_51_473 ();
 decap_12 FILLER_51_485 ();
 fill_4 FILLER_51_497 ();
 fill_2 FILLER_51_501 ();
 fill_1 FILLER_51_503 ();
 decap_12 FILLER_51_505 ();
 decap_12 FILLER_51_517 ();
 decap_12 FILLER_51_529 ();
 decap_12 FILLER_51_541 ();
 fill_4 FILLER_51_553 ();
 fill_2 FILLER_51_557 ();
 fill_1 FILLER_51_559 ();
 decap_12 FILLER_51_561 ();
 decap_12 FILLER_51_573 ();
 decap_12 FILLER_51_585 ();
 decap_12 FILLER_51_597 ();
 fill_4 FILLER_51_609 ();
 fill_2 FILLER_51_613 ();
 fill_1 FILLER_51_615 ();
 fill_4 FILLER_51_617 ();
 decap_12 FILLER_52_3 ();
 decap_12 FILLER_52_15 ();
 fill_1 FILLER_52_27 ();
 decap_12 FILLER_52_29 ();
 decap_12 FILLER_52_41 ();
 decap_12 FILLER_52_53 ();
 decap_12 FILLER_52_65 ();
 fill_4 FILLER_52_77 ();
 fill_2 FILLER_52_81 ();
 fill_1 FILLER_52_83 ();
 decap_12 FILLER_52_85 ();
 decap_12 FILLER_52_97 ();
 decap_12 FILLER_52_109 ();
 decap_12 FILLER_52_121 ();
 fill_4 FILLER_52_133 ();
 fill_2 FILLER_52_137 ();
 fill_1 FILLER_52_139 ();
 decap_12 FILLER_52_141 ();
 decap_12 FILLER_52_153 ();
 decap_12 FILLER_52_165 ();
 decap_12 FILLER_52_177 ();
 fill_4 FILLER_52_189 ();
 fill_2 FILLER_52_193 ();
 fill_1 FILLER_52_195 ();
 decap_12 FILLER_52_197 ();
 decap_12 FILLER_52_209 ();
 decap_12 FILLER_52_221 ();
 decap_12 FILLER_52_233 ();
 fill_4 FILLER_52_245 ();
 fill_2 FILLER_52_249 ();
 fill_1 FILLER_52_251 ();
 decap_12 FILLER_52_253 ();
 decap_12 FILLER_52_265 ();
 decap_12 FILLER_52_277 ();
 decap_12 FILLER_52_289 ();
 fill_4 FILLER_52_301 ();
 fill_2 FILLER_52_305 ();
 fill_1 FILLER_52_307 ();
 decap_12 FILLER_52_309 ();
 decap_12 FILLER_52_321 ();
 decap_12 FILLER_52_333 ();
 decap_12 FILLER_52_345 ();
 fill_4 FILLER_52_357 ();
 fill_2 FILLER_52_361 ();
 fill_1 FILLER_52_363 ();
 decap_12 FILLER_52_365 ();
 decap_12 FILLER_52_377 ();
 decap_12 FILLER_52_389 ();
 decap_12 FILLER_52_401 ();
 fill_4 FILLER_52_413 ();
 fill_2 FILLER_52_417 ();
 fill_1 FILLER_52_419 ();
 decap_12 FILLER_52_421 ();
 decap_12 FILLER_52_433 ();
 decap_12 FILLER_52_445 ();
 decap_12 FILLER_52_457 ();
 fill_4 FILLER_52_469 ();
 fill_2 FILLER_52_473 ();
 fill_1 FILLER_52_475 ();
 decap_12 FILLER_52_477 ();
 decap_12 FILLER_52_489 ();
 decap_12 FILLER_52_501 ();
 decap_12 FILLER_52_513 ();
 fill_4 FILLER_52_525 ();
 fill_2 FILLER_52_529 ();
 fill_1 FILLER_52_531 ();
 decap_12 FILLER_52_533 ();
 decap_12 FILLER_52_545 ();
 decap_12 FILLER_52_557 ();
 decap_12 FILLER_52_569 ();
 fill_4 FILLER_52_581 ();
 fill_2 FILLER_52_585 ();
 fill_1 FILLER_52_587 ();
 decap_12 FILLER_52_589 ();
 decap_12 FILLER_52_601 ();
 decap_12 FILLER_52_613 ();
 decap_12 FILLER_53_3 ();
 decap_12 FILLER_53_15 ();
 decap_12 FILLER_53_27 ();
 decap_12 FILLER_53_39 ();
 fill_4 FILLER_53_51 ();
 fill_1 FILLER_53_55 ();
 decap_12 FILLER_53_57 ();
 decap_12 FILLER_53_69 ();
 decap_12 FILLER_53_81 ();
 decap_12 FILLER_53_93 ();
 fill_4 FILLER_53_105 ();
 fill_2 FILLER_53_109 ();
 fill_1 FILLER_53_111 ();
 decap_12 FILLER_53_113 ();
 decap_12 FILLER_53_125 ();
 decap_12 FILLER_53_137 ();
 decap_12 FILLER_53_149 ();
 fill_4 FILLER_53_161 ();
 fill_2 FILLER_53_165 ();
 fill_1 FILLER_53_167 ();
 decap_12 FILLER_53_169 ();
 decap_12 FILLER_53_181 ();
 decap_12 FILLER_53_193 ();
 decap_12 FILLER_53_205 ();
 fill_4 FILLER_53_217 ();
 fill_2 FILLER_53_221 ();
 fill_1 FILLER_53_223 ();
 decap_12 FILLER_53_225 ();
 decap_12 FILLER_53_237 ();
 decap_12 FILLER_53_249 ();
 decap_12 FILLER_53_261 ();
 fill_4 FILLER_53_273 ();
 fill_2 FILLER_53_277 ();
 fill_1 FILLER_53_279 ();
 decap_12 FILLER_53_281 ();
 decap_12 FILLER_53_293 ();
 decap_12 FILLER_53_305 ();
 decap_12 FILLER_53_317 ();
 fill_4 FILLER_53_329 ();
 fill_2 FILLER_53_333 ();
 fill_1 FILLER_53_335 ();
 decap_12 FILLER_53_337 ();
 decap_12 FILLER_53_349 ();
 decap_12 FILLER_53_361 ();
 decap_12 FILLER_53_373 ();
 fill_4 FILLER_53_385 ();
 fill_2 FILLER_53_389 ();
 fill_1 FILLER_53_391 ();
 decap_12 FILLER_53_393 ();
 decap_12 FILLER_53_405 ();
 decap_12 FILLER_53_417 ();
 decap_12 FILLER_53_429 ();
 fill_4 FILLER_53_441 ();
 fill_2 FILLER_53_445 ();
 fill_1 FILLER_53_447 ();
 decap_12 FILLER_53_449 ();
 decap_12 FILLER_53_461 ();
 decap_12 FILLER_53_473 ();
 decap_12 FILLER_53_485 ();
 fill_4 FILLER_53_497 ();
 fill_2 FILLER_53_501 ();
 fill_1 FILLER_53_503 ();
 decap_12 FILLER_53_505 ();
 decap_12 FILLER_53_517 ();
 decap_12 FILLER_53_529 ();
 decap_12 FILLER_53_541 ();
 fill_4 FILLER_53_553 ();
 fill_2 FILLER_53_557 ();
 fill_1 FILLER_53_559 ();
 decap_12 FILLER_53_561 ();
 decap_12 FILLER_53_573 ();
 decap_12 FILLER_53_585 ();
 decap_12 FILLER_53_597 ();
 fill_4 FILLER_53_609 ();
 fill_2 FILLER_53_613 ();
 fill_1 FILLER_53_615 ();
 fill_8 FILLER_53_617 ();
 decap_12 FILLER_54_3 ();
 decap_12 FILLER_54_15 ();
 fill_1 FILLER_54_27 ();
 decap_12 FILLER_54_29 ();
 decap_12 FILLER_54_41 ();
 decap_12 FILLER_54_53 ();
 decap_12 FILLER_54_65 ();
 fill_4 FILLER_54_77 ();
 fill_2 FILLER_54_81 ();
 fill_1 FILLER_54_83 ();
 decap_12 FILLER_54_85 ();
 decap_12 FILLER_54_97 ();
 decap_12 FILLER_54_109 ();
 decap_12 FILLER_54_121 ();
 fill_4 FILLER_54_133 ();
 fill_2 FILLER_54_137 ();
 fill_1 FILLER_54_139 ();
 decap_12 FILLER_54_141 ();
 decap_12 FILLER_54_153 ();
 decap_12 FILLER_54_165 ();
 decap_12 FILLER_54_177 ();
 fill_4 FILLER_54_189 ();
 fill_2 FILLER_54_193 ();
 fill_1 FILLER_54_195 ();
 decap_12 FILLER_54_197 ();
 decap_12 FILLER_54_209 ();
 decap_12 FILLER_54_221 ();
 decap_12 FILLER_54_233 ();
 fill_4 FILLER_54_245 ();
 fill_2 FILLER_54_249 ();
 fill_1 FILLER_54_251 ();
 decap_12 FILLER_54_253 ();
 decap_12 FILLER_54_265 ();
 decap_12 FILLER_54_277 ();
 decap_12 FILLER_54_289 ();
 fill_4 FILLER_54_301 ();
 fill_2 FILLER_54_305 ();
 fill_1 FILLER_54_307 ();
 decap_12 FILLER_54_309 ();
 decap_12 FILLER_54_321 ();
 decap_12 FILLER_54_333 ();
 decap_12 FILLER_54_345 ();
 fill_4 FILLER_54_357 ();
 fill_2 FILLER_54_361 ();
 fill_1 FILLER_54_363 ();
 decap_12 FILLER_54_365 ();
 decap_12 FILLER_54_377 ();
 decap_12 FILLER_54_389 ();
 decap_12 FILLER_54_401 ();
 fill_4 FILLER_54_413 ();
 fill_2 FILLER_54_417 ();
 fill_1 FILLER_54_419 ();
 decap_12 FILLER_54_421 ();
 decap_12 FILLER_54_433 ();
 decap_12 FILLER_54_445 ();
 decap_12 FILLER_54_457 ();
 fill_4 FILLER_54_469 ();
 fill_2 FILLER_54_473 ();
 fill_1 FILLER_54_475 ();
 decap_12 FILLER_54_477 ();
 decap_12 FILLER_54_489 ();
 decap_12 FILLER_54_501 ();
 decap_12 FILLER_54_513 ();
 fill_4 FILLER_54_525 ();
 fill_2 FILLER_54_529 ();
 fill_1 FILLER_54_531 ();
 decap_12 FILLER_54_533 ();
 decap_12 FILLER_54_545 ();
 decap_12 FILLER_54_557 ();
 decap_12 FILLER_54_569 ();
 fill_4 FILLER_54_581 ();
 fill_2 FILLER_54_585 ();
 fill_1 FILLER_54_587 ();
 decap_12 FILLER_54_589 ();
 decap_12 FILLER_54_601 ();
 decap_12 FILLER_54_613 ();
 decap_12 FILLER_55_3 ();
 decap_12 FILLER_55_15 ();
 decap_12 FILLER_55_27 ();
 decap_12 FILLER_55_39 ();
 fill_4 FILLER_55_51 ();
 fill_1 FILLER_55_55 ();
 decap_12 FILLER_55_57 ();
 decap_12 FILLER_55_69 ();
 decap_12 FILLER_55_81 ();
 decap_12 FILLER_55_93 ();
 fill_4 FILLER_55_105 ();
 fill_2 FILLER_55_109 ();
 fill_1 FILLER_55_111 ();
 decap_12 FILLER_55_113 ();
 decap_12 FILLER_55_125 ();
 decap_12 FILLER_55_137 ();
 decap_12 FILLER_55_149 ();
 fill_4 FILLER_55_161 ();
 fill_2 FILLER_55_165 ();
 fill_1 FILLER_55_167 ();
 decap_12 FILLER_55_169 ();
 decap_12 FILLER_55_181 ();
 decap_12 FILLER_55_193 ();
 decap_12 FILLER_55_205 ();
 fill_4 FILLER_55_217 ();
 fill_2 FILLER_55_221 ();
 fill_1 FILLER_55_223 ();
 decap_12 FILLER_55_225 ();
 decap_12 FILLER_55_237 ();
 decap_12 FILLER_55_249 ();
 decap_12 FILLER_55_261 ();
 fill_4 FILLER_55_273 ();
 fill_2 FILLER_55_277 ();
 fill_1 FILLER_55_279 ();
 decap_12 FILLER_55_281 ();
 decap_12 FILLER_55_293 ();
 decap_12 FILLER_55_305 ();
 decap_12 FILLER_55_317 ();
 fill_4 FILLER_55_329 ();
 fill_2 FILLER_55_333 ();
 fill_1 FILLER_55_335 ();
 decap_12 FILLER_55_337 ();
 decap_12 FILLER_55_349 ();
 decap_12 FILLER_55_361 ();
 decap_12 FILLER_55_373 ();
 fill_4 FILLER_55_385 ();
 fill_2 FILLER_55_389 ();
 fill_1 FILLER_55_391 ();
 decap_12 FILLER_55_393 ();
 decap_12 FILLER_55_405 ();
 decap_12 FILLER_55_417 ();
 decap_12 FILLER_55_429 ();
 fill_4 FILLER_55_441 ();
 fill_2 FILLER_55_445 ();
 fill_1 FILLER_55_447 ();
 decap_12 FILLER_55_449 ();
 decap_12 FILLER_55_461 ();
 decap_12 FILLER_55_473 ();
 decap_12 FILLER_55_485 ();
 fill_4 FILLER_55_497 ();
 fill_2 FILLER_55_501 ();
 fill_1 FILLER_55_503 ();
 decap_12 FILLER_55_505 ();
 decap_12 FILLER_55_517 ();
 decap_12 FILLER_55_529 ();
 decap_12 FILLER_55_541 ();
 fill_4 FILLER_55_553 ();
 fill_2 FILLER_55_557 ();
 fill_1 FILLER_55_559 ();
 decap_12 FILLER_55_561 ();
 decap_12 FILLER_55_573 ();
 decap_12 FILLER_55_585 ();
 decap_12 FILLER_55_597 ();
 fill_4 FILLER_55_609 ();
 fill_2 FILLER_55_613 ();
 fill_1 FILLER_55_615 ();
 fill_8 FILLER_55_617 ();
 decap_12 FILLER_56_3 ();
 decap_12 FILLER_56_15 ();
 fill_1 FILLER_56_27 ();
 decap_12 FILLER_56_29 ();
 decap_12 FILLER_56_41 ();
 decap_12 FILLER_56_53 ();
 decap_12 FILLER_56_65 ();
 fill_4 FILLER_56_77 ();
 fill_2 FILLER_56_81 ();
 fill_1 FILLER_56_83 ();
 decap_12 FILLER_56_85 ();
 decap_12 FILLER_56_97 ();
 decap_12 FILLER_56_109 ();
 decap_12 FILLER_56_121 ();
 fill_4 FILLER_56_133 ();
 fill_2 FILLER_56_137 ();
 fill_1 FILLER_56_139 ();
 decap_12 FILLER_56_141 ();
 decap_12 FILLER_56_153 ();
 decap_12 FILLER_56_165 ();
 decap_12 FILLER_56_177 ();
 fill_4 FILLER_56_189 ();
 fill_2 FILLER_56_193 ();
 fill_1 FILLER_56_195 ();
 decap_12 FILLER_56_197 ();
 decap_12 FILLER_56_209 ();
 decap_12 FILLER_56_221 ();
 decap_12 FILLER_56_233 ();
 fill_4 FILLER_56_245 ();
 fill_2 FILLER_56_249 ();
 fill_1 FILLER_56_251 ();
 decap_12 FILLER_56_253 ();
 decap_12 FILLER_56_265 ();
 decap_12 FILLER_56_277 ();
 decap_12 FILLER_56_289 ();
 fill_4 FILLER_56_301 ();
 fill_2 FILLER_56_305 ();
 fill_1 FILLER_56_307 ();
 decap_12 FILLER_56_309 ();
 decap_12 FILLER_56_321 ();
 decap_12 FILLER_56_333 ();
 decap_12 FILLER_56_345 ();
 fill_4 FILLER_56_357 ();
 fill_2 FILLER_56_361 ();
 fill_1 FILLER_56_363 ();
 decap_12 FILLER_56_365 ();
 decap_12 FILLER_56_377 ();
 decap_12 FILLER_56_389 ();
 decap_12 FILLER_56_401 ();
 fill_4 FILLER_56_413 ();
 fill_2 FILLER_56_417 ();
 fill_1 FILLER_56_419 ();
 decap_12 FILLER_56_421 ();
 decap_12 FILLER_56_433 ();
 decap_12 FILLER_56_445 ();
 decap_12 FILLER_56_457 ();
 fill_4 FILLER_56_469 ();
 fill_2 FILLER_56_473 ();
 fill_1 FILLER_56_475 ();
 decap_12 FILLER_56_477 ();
 decap_12 FILLER_56_489 ();
 decap_12 FILLER_56_501 ();
 decap_12 FILLER_56_513 ();
 fill_4 FILLER_56_525 ();
 fill_2 FILLER_56_529 ();
 fill_1 FILLER_56_531 ();
 decap_12 FILLER_56_533 ();
 decap_12 FILLER_56_545 ();
 decap_12 FILLER_56_557 ();
 decap_12 FILLER_56_569 ();
 fill_4 FILLER_56_581 ();
 fill_2 FILLER_56_585 ();
 fill_1 FILLER_56_587 ();
 decap_12 FILLER_56_589 ();
 decap_12 FILLER_56_601 ();
 decap_12 FILLER_56_613 ();
 decap_12 FILLER_57_3 ();
 decap_12 FILLER_57_15 ();
 decap_12 FILLER_57_27 ();
 decap_12 FILLER_57_39 ();
 fill_4 FILLER_57_51 ();
 fill_1 FILLER_57_55 ();
 decap_12 FILLER_57_57 ();
 decap_12 FILLER_57_69 ();
 decap_12 FILLER_57_81 ();
 decap_12 FILLER_57_93 ();
 fill_4 FILLER_57_105 ();
 fill_2 FILLER_57_109 ();
 fill_1 FILLER_57_111 ();
 decap_12 FILLER_57_113 ();
 decap_12 FILLER_57_125 ();
 decap_12 FILLER_57_137 ();
 decap_12 FILLER_57_149 ();
 fill_4 FILLER_57_161 ();
 fill_2 FILLER_57_165 ();
 fill_1 FILLER_57_167 ();
 decap_12 FILLER_57_169 ();
 decap_12 FILLER_57_181 ();
 decap_12 FILLER_57_193 ();
 decap_12 FILLER_57_205 ();
 fill_4 FILLER_57_217 ();
 fill_2 FILLER_57_221 ();
 fill_1 FILLER_57_223 ();
 decap_12 FILLER_57_225 ();
 decap_12 FILLER_57_237 ();
 decap_12 FILLER_57_249 ();
 decap_12 FILLER_57_261 ();
 fill_4 FILLER_57_273 ();
 fill_2 FILLER_57_277 ();
 fill_1 FILLER_57_279 ();
 decap_12 FILLER_57_281 ();
 decap_12 FILLER_57_293 ();
 decap_12 FILLER_57_305 ();
 decap_12 FILLER_57_317 ();
 fill_4 FILLER_57_329 ();
 fill_2 FILLER_57_333 ();
 fill_1 FILLER_57_335 ();
 decap_12 FILLER_57_337 ();
 decap_12 FILLER_57_349 ();
 decap_12 FILLER_57_361 ();
 decap_12 FILLER_57_373 ();
 fill_4 FILLER_57_385 ();
 fill_2 FILLER_57_389 ();
 fill_1 FILLER_57_391 ();
 decap_12 FILLER_57_393 ();
 decap_12 FILLER_57_405 ();
 decap_12 FILLER_57_417 ();
 decap_12 FILLER_57_429 ();
 fill_4 FILLER_57_441 ();
 fill_2 FILLER_57_445 ();
 fill_1 FILLER_57_447 ();
 decap_12 FILLER_57_449 ();
 decap_12 FILLER_57_461 ();
 decap_12 FILLER_57_473 ();
 decap_12 FILLER_57_485 ();
 fill_4 FILLER_57_497 ();
 fill_2 FILLER_57_501 ();
 fill_1 FILLER_57_503 ();
 decap_12 FILLER_57_505 ();
 decap_12 FILLER_57_517 ();
 decap_12 FILLER_57_529 ();
 decap_12 FILLER_57_541 ();
 fill_4 FILLER_57_553 ();
 fill_2 FILLER_57_557 ();
 fill_1 FILLER_57_559 ();
 decap_12 FILLER_57_561 ();
 decap_12 FILLER_57_573 ();
 decap_12 FILLER_57_585 ();
 decap_12 FILLER_57_597 ();
 fill_4 FILLER_57_609 ();
 fill_2 FILLER_57_613 ();
 fill_1 FILLER_57_615 ();
 fill_8 FILLER_57_617 ();
 decap_12 FILLER_58_3 ();
 decap_12 FILLER_58_15 ();
 fill_1 FILLER_58_27 ();
 decap_12 FILLER_58_29 ();
 decap_12 FILLER_58_41 ();
 decap_12 FILLER_58_53 ();
 decap_12 FILLER_58_65 ();
 fill_4 FILLER_58_77 ();
 fill_2 FILLER_58_81 ();
 fill_1 FILLER_58_83 ();
 decap_12 FILLER_58_85 ();
 decap_12 FILLER_58_97 ();
 decap_12 FILLER_58_109 ();
 decap_12 FILLER_58_121 ();
 fill_4 FILLER_58_133 ();
 fill_2 FILLER_58_137 ();
 fill_1 FILLER_58_139 ();
 decap_12 FILLER_58_141 ();
 decap_12 FILLER_58_153 ();
 decap_12 FILLER_58_165 ();
 decap_12 FILLER_58_177 ();
 fill_4 FILLER_58_189 ();
 fill_2 FILLER_58_193 ();
 fill_1 FILLER_58_195 ();
 decap_12 FILLER_58_197 ();
 decap_12 FILLER_58_209 ();
 decap_12 FILLER_58_221 ();
 decap_12 FILLER_58_233 ();
 fill_4 FILLER_58_245 ();
 fill_2 FILLER_58_249 ();
 fill_1 FILLER_58_251 ();
 decap_12 FILLER_58_253 ();
 decap_12 FILLER_58_265 ();
 decap_12 FILLER_58_277 ();
 decap_12 FILLER_58_289 ();
 fill_4 FILLER_58_301 ();
 fill_2 FILLER_58_305 ();
 fill_1 FILLER_58_307 ();
 decap_12 FILLER_58_309 ();
 decap_12 FILLER_58_321 ();
 decap_12 FILLER_58_333 ();
 decap_12 FILLER_58_345 ();
 fill_4 FILLER_58_357 ();
 fill_2 FILLER_58_361 ();
 fill_1 FILLER_58_363 ();
 decap_12 FILLER_58_365 ();
 decap_12 FILLER_58_377 ();
 decap_12 FILLER_58_389 ();
 decap_12 FILLER_58_401 ();
 fill_4 FILLER_58_413 ();
 fill_2 FILLER_58_417 ();
 fill_1 FILLER_58_419 ();
 decap_12 FILLER_58_421 ();
 decap_12 FILLER_58_433 ();
 decap_12 FILLER_58_445 ();
 decap_12 FILLER_58_457 ();
 fill_4 FILLER_58_469 ();
 fill_2 FILLER_58_473 ();
 fill_1 FILLER_58_475 ();
 decap_12 FILLER_58_477 ();
 decap_12 FILLER_58_489 ();
 decap_12 FILLER_58_501 ();
 decap_12 FILLER_58_513 ();
 fill_4 FILLER_58_525 ();
 fill_2 FILLER_58_529 ();
 fill_1 FILLER_58_531 ();
 decap_12 FILLER_58_533 ();
 decap_12 FILLER_58_545 ();
 decap_12 FILLER_58_557 ();
 decap_12 FILLER_58_569 ();
 fill_4 FILLER_58_581 ();
 fill_2 FILLER_58_585 ();
 fill_1 FILLER_58_587 ();
 decap_12 FILLER_58_589 ();
 decap_12 FILLER_58_601 ();
 decap_12 FILLER_58_613 ();
 decap_12 FILLER_59_3 ();
 decap_12 FILLER_59_15 ();
 decap_12 FILLER_59_27 ();
 decap_12 FILLER_59_39 ();
 fill_4 FILLER_59_51 ();
 fill_1 FILLER_59_55 ();
 decap_12 FILLER_59_57 ();
 decap_12 FILLER_59_69 ();
 decap_12 FILLER_59_81 ();
 decap_12 FILLER_59_93 ();
 fill_4 FILLER_59_105 ();
 fill_2 FILLER_59_109 ();
 fill_1 FILLER_59_111 ();
 decap_12 FILLER_59_113 ();
 decap_12 FILLER_59_125 ();
 decap_12 FILLER_59_137 ();
 decap_12 FILLER_59_149 ();
 fill_4 FILLER_59_161 ();
 fill_2 FILLER_59_165 ();
 fill_1 FILLER_59_167 ();
 decap_12 FILLER_59_169 ();
 decap_12 FILLER_59_181 ();
 decap_12 FILLER_59_193 ();
 decap_12 FILLER_59_205 ();
 fill_4 FILLER_59_217 ();
 fill_2 FILLER_59_221 ();
 fill_1 FILLER_59_223 ();
 decap_12 FILLER_59_225 ();
 decap_12 FILLER_59_237 ();
 decap_12 FILLER_59_249 ();
 decap_12 FILLER_59_261 ();
 fill_4 FILLER_59_273 ();
 fill_2 FILLER_59_277 ();
 fill_1 FILLER_59_279 ();
 decap_12 FILLER_59_281 ();
 decap_12 FILLER_59_293 ();
 decap_12 FILLER_59_305 ();
 decap_12 FILLER_59_317 ();
 fill_4 FILLER_59_329 ();
 fill_2 FILLER_59_333 ();
 fill_1 FILLER_59_335 ();
 decap_12 FILLER_59_337 ();
 decap_12 FILLER_59_349 ();
 decap_12 FILLER_59_361 ();
 decap_12 FILLER_59_373 ();
 fill_4 FILLER_59_385 ();
 fill_2 FILLER_59_389 ();
 fill_1 FILLER_59_391 ();
 decap_12 FILLER_59_393 ();
 decap_12 FILLER_59_405 ();
 decap_12 FILLER_59_417 ();
 decap_12 FILLER_59_429 ();
 fill_4 FILLER_59_441 ();
 fill_2 FILLER_59_445 ();
 fill_1 FILLER_59_447 ();
 decap_12 FILLER_59_449 ();
 decap_12 FILLER_59_461 ();
 decap_12 FILLER_59_473 ();
 decap_12 FILLER_59_485 ();
 fill_4 FILLER_59_497 ();
 fill_2 FILLER_59_501 ();
 fill_1 FILLER_59_503 ();
 decap_12 FILLER_59_505 ();
 decap_12 FILLER_59_517 ();
 decap_12 FILLER_59_529 ();
 decap_12 FILLER_59_541 ();
 fill_4 FILLER_59_553 ();
 fill_2 FILLER_59_557 ();
 fill_1 FILLER_59_559 ();
 decap_12 FILLER_59_561 ();
 decap_12 FILLER_59_573 ();
 decap_12 FILLER_59_585 ();
 decap_12 FILLER_59_597 ();
 fill_4 FILLER_59_609 ();
 fill_2 FILLER_59_613 ();
 fill_1 FILLER_59_615 ();
 fill_8 FILLER_59_617 ();
 decap_12 FILLER_60_3 ();
 decap_12 FILLER_60_15 ();
 fill_1 FILLER_60_27 ();
 decap_12 FILLER_60_29 ();
 decap_12 FILLER_60_41 ();
 decap_12 FILLER_60_53 ();
 decap_12 FILLER_60_65 ();
 fill_4 FILLER_60_77 ();
 fill_2 FILLER_60_81 ();
 fill_1 FILLER_60_83 ();
 decap_12 FILLER_60_85 ();
 decap_12 FILLER_60_97 ();
 decap_12 FILLER_60_109 ();
 decap_12 FILLER_60_121 ();
 fill_4 FILLER_60_133 ();
 fill_2 FILLER_60_137 ();
 fill_1 FILLER_60_139 ();
 decap_12 FILLER_60_141 ();
 decap_12 FILLER_60_153 ();
 decap_12 FILLER_60_165 ();
 decap_12 FILLER_60_177 ();
 fill_4 FILLER_60_189 ();
 fill_2 FILLER_60_193 ();
 fill_1 FILLER_60_195 ();
 decap_12 FILLER_60_197 ();
 decap_12 FILLER_60_209 ();
 decap_12 FILLER_60_221 ();
 decap_12 FILLER_60_233 ();
 fill_4 FILLER_60_245 ();
 fill_2 FILLER_60_249 ();
 fill_1 FILLER_60_251 ();
 decap_12 FILLER_60_253 ();
 decap_12 FILLER_60_265 ();
 decap_12 FILLER_60_277 ();
 decap_12 FILLER_60_289 ();
 fill_4 FILLER_60_301 ();
 fill_2 FILLER_60_305 ();
 fill_1 FILLER_60_307 ();
 decap_12 FILLER_60_309 ();
 decap_12 FILLER_60_321 ();
 decap_12 FILLER_60_333 ();
 decap_12 FILLER_60_345 ();
 fill_4 FILLER_60_357 ();
 fill_2 FILLER_60_361 ();
 fill_1 FILLER_60_363 ();
 decap_12 FILLER_60_365 ();
 decap_12 FILLER_60_377 ();
 decap_12 FILLER_60_389 ();
 decap_12 FILLER_60_401 ();
 fill_4 FILLER_60_413 ();
 fill_2 FILLER_60_417 ();
 fill_1 FILLER_60_419 ();
 decap_12 FILLER_60_421 ();
 decap_12 FILLER_60_433 ();
 decap_12 FILLER_60_445 ();
 decap_12 FILLER_60_457 ();
 fill_4 FILLER_60_469 ();
 fill_2 FILLER_60_473 ();
 fill_1 FILLER_60_475 ();
 decap_12 FILLER_60_477 ();
 decap_12 FILLER_60_489 ();
 decap_12 FILLER_60_501 ();
 decap_12 FILLER_60_513 ();
 fill_4 FILLER_60_525 ();
 fill_2 FILLER_60_529 ();
 fill_1 FILLER_60_531 ();
 decap_12 FILLER_60_533 ();
 decap_12 FILLER_60_545 ();
 decap_12 FILLER_60_557 ();
 decap_12 FILLER_60_569 ();
 fill_4 FILLER_60_581 ();
 fill_2 FILLER_60_585 ();
 fill_1 FILLER_60_587 ();
 decap_12 FILLER_60_589 ();
 decap_12 FILLER_60_601 ();
 decap_12 FILLER_60_613 ();
 decap_12 FILLER_61_3 ();
 decap_12 FILLER_61_15 ();
 decap_12 FILLER_61_27 ();
 decap_12 FILLER_61_39 ();
 fill_4 FILLER_61_51 ();
 fill_1 FILLER_61_55 ();
 decap_12 FILLER_61_57 ();
 decap_12 FILLER_61_69 ();
 decap_12 FILLER_61_81 ();
 decap_12 FILLER_61_93 ();
 fill_4 FILLER_61_105 ();
 fill_2 FILLER_61_109 ();
 fill_1 FILLER_61_111 ();
 decap_12 FILLER_61_113 ();
 decap_12 FILLER_61_125 ();
 decap_12 FILLER_61_137 ();
 decap_12 FILLER_61_149 ();
 fill_4 FILLER_61_161 ();
 fill_2 FILLER_61_165 ();
 fill_1 FILLER_61_167 ();
 decap_12 FILLER_61_169 ();
 decap_12 FILLER_61_181 ();
 decap_12 FILLER_61_193 ();
 decap_12 FILLER_61_205 ();
 fill_4 FILLER_61_217 ();
 fill_2 FILLER_61_221 ();
 fill_1 FILLER_61_223 ();
 decap_12 FILLER_61_225 ();
 decap_12 FILLER_61_237 ();
 decap_12 FILLER_61_249 ();
 decap_12 FILLER_61_261 ();
 fill_4 FILLER_61_273 ();
 fill_2 FILLER_61_277 ();
 fill_1 FILLER_61_279 ();
 decap_12 FILLER_61_281 ();
 decap_12 FILLER_61_293 ();
 decap_12 FILLER_61_305 ();
 decap_12 FILLER_61_317 ();
 fill_4 FILLER_61_329 ();
 fill_2 FILLER_61_333 ();
 fill_1 FILLER_61_335 ();
 decap_12 FILLER_61_337 ();
 decap_12 FILLER_61_349 ();
 decap_12 FILLER_61_361 ();
 decap_12 FILLER_61_373 ();
 fill_4 FILLER_61_385 ();
 fill_2 FILLER_61_389 ();
 fill_1 FILLER_61_391 ();
 decap_12 FILLER_61_393 ();
 decap_12 FILLER_61_405 ();
 decap_12 FILLER_61_417 ();
 decap_12 FILLER_61_429 ();
 fill_4 FILLER_61_441 ();
 fill_2 FILLER_61_445 ();
 fill_1 FILLER_61_447 ();
 decap_12 FILLER_61_449 ();
 decap_12 FILLER_61_461 ();
 decap_12 FILLER_61_473 ();
 decap_12 FILLER_61_485 ();
 fill_4 FILLER_61_497 ();
 fill_2 FILLER_61_501 ();
 fill_1 FILLER_61_503 ();
 decap_12 FILLER_61_505 ();
 decap_12 FILLER_61_517 ();
 decap_12 FILLER_61_529 ();
 decap_12 FILLER_61_541 ();
 fill_4 FILLER_61_553 ();
 fill_2 FILLER_61_557 ();
 fill_1 FILLER_61_559 ();
 decap_12 FILLER_61_561 ();
 decap_12 FILLER_61_573 ();
 decap_12 FILLER_61_585 ();
 decap_12 FILLER_61_597 ();
 fill_4 FILLER_61_609 ();
 fill_2 FILLER_61_613 ();
 fill_1 FILLER_61_615 ();
 fill_8 FILLER_61_617 ();
 decap_12 FILLER_62_3 ();
 decap_12 FILLER_62_15 ();
 fill_1 FILLER_62_27 ();
 decap_12 FILLER_62_29 ();
 decap_12 FILLER_62_41 ();
 decap_12 FILLER_62_53 ();
 decap_12 FILLER_62_65 ();
 fill_4 FILLER_62_77 ();
 fill_2 FILLER_62_81 ();
 fill_1 FILLER_62_83 ();
 decap_12 FILLER_62_85 ();
 decap_12 FILLER_62_97 ();
 decap_12 FILLER_62_109 ();
 decap_12 FILLER_62_121 ();
 fill_4 FILLER_62_133 ();
 fill_2 FILLER_62_137 ();
 fill_1 FILLER_62_139 ();
 decap_12 FILLER_62_141 ();
 decap_12 FILLER_62_153 ();
 decap_12 FILLER_62_165 ();
 decap_12 FILLER_62_177 ();
 fill_4 FILLER_62_189 ();
 fill_2 FILLER_62_193 ();
 fill_1 FILLER_62_195 ();
 decap_12 FILLER_62_197 ();
 decap_12 FILLER_62_209 ();
 decap_12 FILLER_62_221 ();
 decap_12 FILLER_62_233 ();
 fill_4 FILLER_62_245 ();
 fill_2 FILLER_62_249 ();
 fill_1 FILLER_62_251 ();
 decap_12 FILLER_62_253 ();
 decap_12 FILLER_62_265 ();
 decap_12 FILLER_62_277 ();
 decap_12 FILLER_62_289 ();
 fill_4 FILLER_62_301 ();
 fill_2 FILLER_62_305 ();
 fill_1 FILLER_62_307 ();
 decap_12 FILLER_62_309 ();
 decap_12 FILLER_62_321 ();
 decap_12 FILLER_62_333 ();
 decap_12 FILLER_62_345 ();
 fill_4 FILLER_62_357 ();
 fill_2 FILLER_62_361 ();
 fill_1 FILLER_62_363 ();
 decap_12 FILLER_62_365 ();
 decap_12 FILLER_62_377 ();
 decap_12 FILLER_62_389 ();
 decap_12 FILLER_62_401 ();
 fill_4 FILLER_62_413 ();
 fill_2 FILLER_62_417 ();
 fill_1 FILLER_62_419 ();
 decap_12 FILLER_62_421 ();
 decap_12 FILLER_62_433 ();
 decap_12 FILLER_62_445 ();
 decap_12 FILLER_62_457 ();
 fill_4 FILLER_62_469 ();
 fill_2 FILLER_62_473 ();
 fill_1 FILLER_62_475 ();
 decap_12 FILLER_62_477 ();
 decap_12 FILLER_62_489 ();
 decap_12 FILLER_62_501 ();
 decap_12 FILLER_62_513 ();
 fill_4 FILLER_62_525 ();
 fill_2 FILLER_62_529 ();
 fill_1 FILLER_62_531 ();
 decap_12 FILLER_62_533 ();
 decap_12 FILLER_62_545 ();
 decap_12 FILLER_62_557 ();
 decap_12 FILLER_62_569 ();
 fill_4 FILLER_62_581 ();
 fill_2 FILLER_62_585 ();
 fill_1 FILLER_62_587 ();
 decap_12 FILLER_62_589 ();
 decap_12 FILLER_62_601 ();
 decap_12 FILLER_62_613 ();
 decap_12 FILLER_63_3 ();
 decap_12 FILLER_63_15 ();
 decap_12 FILLER_63_27 ();
 decap_12 FILLER_63_39 ();
 fill_4 FILLER_63_51 ();
 fill_1 FILLER_63_55 ();
 decap_12 FILLER_63_57 ();
 decap_12 FILLER_63_69 ();
 decap_12 FILLER_63_81 ();
 decap_12 FILLER_63_93 ();
 fill_4 FILLER_63_105 ();
 fill_2 FILLER_63_109 ();
 fill_1 FILLER_63_111 ();
 decap_12 FILLER_63_113 ();
 decap_12 FILLER_63_125 ();
 decap_12 FILLER_63_137 ();
 decap_12 FILLER_63_149 ();
 fill_4 FILLER_63_161 ();
 fill_2 FILLER_63_165 ();
 fill_1 FILLER_63_167 ();
 decap_12 FILLER_63_169 ();
 decap_12 FILLER_63_181 ();
 decap_12 FILLER_63_193 ();
 decap_12 FILLER_63_205 ();
 fill_4 FILLER_63_217 ();
 fill_2 FILLER_63_221 ();
 fill_1 FILLER_63_223 ();
 decap_12 FILLER_63_225 ();
 decap_12 FILLER_63_237 ();
 decap_12 FILLER_63_249 ();
 decap_12 FILLER_63_261 ();
 fill_4 FILLER_63_273 ();
 fill_2 FILLER_63_277 ();
 fill_1 FILLER_63_279 ();
 decap_12 FILLER_63_281 ();
 decap_12 FILLER_63_293 ();
 decap_12 FILLER_63_305 ();
 decap_12 FILLER_63_317 ();
 fill_4 FILLER_63_329 ();
 fill_2 FILLER_63_333 ();
 fill_1 FILLER_63_335 ();
 decap_12 FILLER_63_337 ();
 decap_12 FILLER_63_349 ();
 decap_12 FILLER_63_361 ();
 decap_12 FILLER_63_373 ();
 fill_4 FILLER_63_385 ();
 fill_2 FILLER_63_389 ();
 fill_1 FILLER_63_391 ();
 decap_12 FILLER_63_393 ();
 decap_12 FILLER_63_405 ();
 decap_12 FILLER_63_417 ();
 decap_12 FILLER_63_429 ();
 fill_4 FILLER_63_441 ();
 fill_2 FILLER_63_445 ();
 fill_1 FILLER_63_447 ();
 decap_12 FILLER_63_449 ();
 decap_12 FILLER_63_461 ();
 decap_12 FILLER_63_473 ();
 decap_12 FILLER_63_485 ();
 fill_4 FILLER_63_497 ();
 fill_2 FILLER_63_501 ();
 fill_1 FILLER_63_503 ();
 decap_12 FILLER_63_505 ();
 decap_12 FILLER_63_517 ();
 decap_12 FILLER_63_529 ();
 decap_12 FILLER_63_541 ();
 fill_4 FILLER_63_553 ();
 fill_2 FILLER_63_557 ();
 fill_1 FILLER_63_559 ();
 decap_12 FILLER_63_561 ();
 decap_12 FILLER_63_573 ();
 decap_12 FILLER_63_585 ();
 decap_12 FILLER_63_597 ();
 fill_4 FILLER_63_609 ();
 fill_2 FILLER_63_613 ();
 fill_1 FILLER_63_615 ();
 fill_8 FILLER_63_617 ();
 decap_12 FILLER_64_3 ();
 decap_12 FILLER_64_15 ();
 fill_1 FILLER_64_27 ();
 decap_12 FILLER_64_29 ();
 decap_12 FILLER_64_41 ();
 decap_12 FILLER_64_53 ();
 decap_12 FILLER_64_65 ();
 fill_4 FILLER_64_77 ();
 fill_2 FILLER_64_81 ();
 fill_1 FILLER_64_83 ();
 decap_12 FILLER_64_85 ();
 decap_12 FILLER_64_97 ();
 decap_12 FILLER_64_109 ();
 decap_12 FILLER_64_121 ();
 fill_4 FILLER_64_133 ();
 fill_2 FILLER_64_137 ();
 fill_1 FILLER_64_139 ();
 decap_12 FILLER_64_141 ();
 decap_12 FILLER_64_153 ();
 decap_12 FILLER_64_165 ();
 decap_12 FILLER_64_177 ();
 fill_4 FILLER_64_189 ();
 fill_2 FILLER_64_193 ();
 fill_1 FILLER_64_195 ();
 decap_12 FILLER_64_197 ();
 decap_12 FILLER_64_209 ();
 decap_12 FILLER_64_221 ();
 decap_12 FILLER_64_233 ();
 fill_4 FILLER_64_245 ();
 fill_2 FILLER_64_249 ();
 fill_1 FILLER_64_251 ();
 decap_12 FILLER_64_253 ();
 decap_12 FILLER_64_265 ();
 decap_12 FILLER_64_277 ();
 decap_12 FILLER_64_289 ();
 fill_4 FILLER_64_301 ();
 fill_2 FILLER_64_305 ();
 fill_1 FILLER_64_307 ();
 decap_12 FILLER_64_309 ();
 decap_12 FILLER_64_321 ();
 decap_12 FILLER_64_333 ();
 decap_12 FILLER_64_345 ();
 fill_4 FILLER_64_357 ();
 fill_2 FILLER_64_361 ();
 fill_1 FILLER_64_363 ();
 decap_12 FILLER_64_365 ();
 decap_12 FILLER_64_377 ();
 decap_12 FILLER_64_389 ();
 decap_12 FILLER_64_401 ();
 fill_4 FILLER_64_413 ();
 fill_2 FILLER_64_417 ();
 fill_1 FILLER_64_419 ();
 decap_12 FILLER_64_421 ();
 decap_12 FILLER_64_433 ();
 decap_12 FILLER_64_445 ();
 decap_12 FILLER_64_457 ();
 fill_4 FILLER_64_469 ();
 fill_2 FILLER_64_473 ();
 fill_1 FILLER_64_475 ();
 decap_12 FILLER_64_477 ();
 decap_12 FILLER_64_489 ();
 decap_12 FILLER_64_501 ();
 decap_12 FILLER_64_513 ();
 fill_4 FILLER_64_525 ();
 fill_2 FILLER_64_529 ();
 fill_1 FILLER_64_531 ();
 decap_12 FILLER_64_533 ();
 decap_12 FILLER_64_545 ();
 decap_12 FILLER_64_557 ();
 decap_12 FILLER_64_569 ();
 fill_4 FILLER_64_581 ();
 fill_2 FILLER_64_585 ();
 fill_1 FILLER_64_587 ();
 decap_12 FILLER_64_589 ();
 decap_12 FILLER_64_601 ();
 decap_12 FILLER_64_613 ();
 decap_12 FILLER_65_3 ();
 decap_12 FILLER_65_15 ();
 decap_12 FILLER_65_27 ();
 decap_12 FILLER_65_39 ();
 fill_4 FILLER_65_51 ();
 fill_1 FILLER_65_55 ();
 decap_12 FILLER_65_57 ();
 decap_12 FILLER_65_69 ();
 decap_12 FILLER_65_81 ();
 decap_12 FILLER_65_93 ();
 fill_4 FILLER_65_105 ();
 fill_2 FILLER_65_109 ();
 fill_1 FILLER_65_111 ();
 decap_12 FILLER_65_113 ();
 decap_12 FILLER_65_125 ();
 decap_12 FILLER_65_137 ();
 decap_12 FILLER_65_149 ();
 fill_4 FILLER_65_161 ();
 fill_2 FILLER_65_165 ();
 fill_1 FILLER_65_167 ();
 decap_12 FILLER_65_169 ();
 decap_12 FILLER_65_181 ();
 decap_12 FILLER_65_193 ();
 decap_12 FILLER_65_205 ();
 fill_4 FILLER_65_217 ();
 fill_2 FILLER_65_221 ();
 fill_1 FILLER_65_223 ();
 decap_12 FILLER_65_225 ();
 decap_12 FILLER_65_237 ();
 decap_12 FILLER_65_249 ();
 decap_12 FILLER_65_261 ();
 fill_4 FILLER_65_273 ();
 fill_2 FILLER_65_277 ();
 fill_1 FILLER_65_279 ();
 decap_12 FILLER_65_281 ();
 decap_12 FILLER_65_293 ();
 decap_12 FILLER_65_305 ();
 decap_12 FILLER_65_317 ();
 fill_4 FILLER_65_329 ();
 fill_2 FILLER_65_333 ();
 fill_1 FILLER_65_335 ();
 decap_12 FILLER_65_337 ();
 decap_12 FILLER_65_349 ();
 decap_12 FILLER_65_361 ();
 decap_12 FILLER_65_373 ();
 fill_4 FILLER_65_385 ();
 fill_2 FILLER_65_389 ();
 fill_1 FILLER_65_391 ();
 decap_12 FILLER_65_393 ();
 decap_12 FILLER_65_405 ();
 decap_12 FILLER_65_417 ();
 decap_12 FILLER_65_429 ();
 fill_4 FILLER_65_441 ();
 fill_2 FILLER_65_445 ();
 fill_1 FILLER_65_447 ();
 decap_12 FILLER_65_449 ();
 decap_12 FILLER_65_461 ();
 decap_12 FILLER_65_473 ();
 decap_12 FILLER_65_485 ();
 fill_4 FILLER_65_497 ();
 fill_2 FILLER_65_501 ();
 fill_1 FILLER_65_503 ();
 decap_12 FILLER_65_505 ();
 decap_12 FILLER_65_517 ();
 decap_12 FILLER_65_529 ();
 decap_12 FILLER_65_541 ();
 fill_4 FILLER_65_553 ();
 fill_2 FILLER_65_557 ();
 fill_1 FILLER_65_559 ();
 decap_12 FILLER_65_561 ();
 decap_12 FILLER_65_573 ();
 decap_12 FILLER_65_585 ();
 decap_12 FILLER_65_597 ();
 fill_4 FILLER_65_609 ();
 fill_2 FILLER_65_613 ();
 fill_1 FILLER_65_615 ();
 fill_8 FILLER_65_617 ();
 decap_12 FILLER_66_3 ();
 decap_12 FILLER_66_15 ();
 fill_1 FILLER_66_27 ();
 decap_12 FILLER_66_29 ();
 decap_12 FILLER_66_41 ();
 decap_12 FILLER_66_53 ();
 decap_12 FILLER_66_65 ();
 fill_4 FILLER_66_77 ();
 fill_2 FILLER_66_81 ();
 fill_1 FILLER_66_83 ();
 decap_12 FILLER_66_85 ();
 decap_12 FILLER_66_97 ();
 decap_12 FILLER_66_109 ();
 decap_12 FILLER_66_121 ();
 fill_4 FILLER_66_133 ();
 fill_2 FILLER_66_137 ();
 fill_1 FILLER_66_139 ();
 decap_12 FILLER_66_141 ();
 decap_12 FILLER_66_153 ();
 decap_12 FILLER_66_165 ();
 decap_12 FILLER_66_177 ();
 fill_4 FILLER_66_189 ();
 fill_2 FILLER_66_193 ();
 fill_1 FILLER_66_195 ();
 decap_12 FILLER_66_197 ();
 decap_12 FILLER_66_209 ();
 decap_12 FILLER_66_221 ();
 decap_12 FILLER_66_233 ();
 fill_4 FILLER_66_245 ();
 fill_2 FILLER_66_249 ();
 fill_1 FILLER_66_251 ();
 decap_12 FILLER_66_253 ();
 decap_12 FILLER_66_265 ();
 decap_12 FILLER_66_277 ();
 decap_12 FILLER_66_289 ();
 fill_4 FILLER_66_301 ();
 fill_2 FILLER_66_305 ();
 fill_1 FILLER_66_307 ();
 decap_12 FILLER_66_309 ();
 decap_12 FILLER_66_321 ();
 decap_12 FILLER_66_333 ();
 decap_12 FILLER_66_345 ();
 fill_4 FILLER_66_357 ();
 fill_2 FILLER_66_361 ();
 fill_1 FILLER_66_363 ();
 decap_12 FILLER_66_365 ();
 decap_12 FILLER_66_377 ();
 decap_12 FILLER_66_389 ();
 decap_12 FILLER_66_401 ();
 fill_4 FILLER_66_413 ();
 fill_2 FILLER_66_417 ();
 fill_1 FILLER_66_419 ();
 decap_12 FILLER_66_421 ();
 decap_12 FILLER_66_433 ();
 decap_12 FILLER_66_445 ();
 decap_12 FILLER_66_457 ();
 fill_4 FILLER_66_469 ();
 fill_2 FILLER_66_473 ();
 fill_1 FILLER_66_475 ();
 decap_12 FILLER_66_477 ();
 decap_12 FILLER_66_489 ();
 decap_12 FILLER_66_501 ();
 decap_12 FILLER_66_513 ();
 fill_4 FILLER_66_525 ();
 fill_2 FILLER_66_529 ();
 fill_1 FILLER_66_531 ();
 decap_12 FILLER_66_533 ();
 decap_12 FILLER_66_545 ();
 decap_12 FILLER_66_557 ();
 decap_12 FILLER_66_569 ();
 fill_4 FILLER_66_581 ();
 fill_2 FILLER_66_585 ();
 fill_1 FILLER_66_587 ();
 decap_12 FILLER_66_589 ();
 decap_12 FILLER_66_601 ();
 decap_12 FILLER_66_613 ();
 decap_12 FILLER_67_3 ();
 decap_12 FILLER_67_15 ();
 decap_12 FILLER_67_27 ();
 decap_12 FILLER_67_39 ();
 fill_4 FILLER_67_51 ();
 fill_1 FILLER_67_55 ();
 decap_12 FILLER_67_57 ();
 decap_12 FILLER_67_69 ();
 decap_12 FILLER_67_81 ();
 decap_12 FILLER_67_93 ();
 fill_4 FILLER_67_105 ();
 fill_2 FILLER_67_109 ();
 fill_1 FILLER_67_111 ();
 decap_12 FILLER_67_113 ();
 decap_12 FILLER_67_125 ();
 decap_12 FILLER_67_137 ();
 decap_12 FILLER_67_149 ();
 fill_4 FILLER_67_161 ();
 fill_2 FILLER_67_165 ();
 fill_1 FILLER_67_167 ();
 decap_12 FILLER_67_169 ();
 decap_12 FILLER_67_181 ();
 decap_12 FILLER_67_193 ();
 decap_12 FILLER_67_205 ();
 fill_4 FILLER_67_217 ();
 fill_2 FILLER_67_221 ();
 fill_1 FILLER_67_223 ();
 decap_12 FILLER_67_225 ();
 decap_12 FILLER_67_237 ();
 decap_12 FILLER_67_249 ();
 decap_12 FILLER_67_261 ();
 fill_4 FILLER_67_273 ();
 fill_2 FILLER_67_277 ();
 fill_1 FILLER_67_279 ();
 decap_12 FILLER_67_281 ();
 decap_12 FILLER_67_293 ();
 decap_12 FILLER_67_305 ();
 decap_12 FILLER_67_317 ();
 fill_4 FILLER_67_329 ();
 fill_2 FILLER_67_333 ();
 fill_1 FILLER_67_335 ();
 decap_12 FILLER_67_337 ();
 decap_12 FILLER_67_349 ();
 decap_12 FILLER_67_361 ();
 decap_12 FILLER_67_373 ();
 fill_4 FILLER_67_385 ();
 fill_2 FILLER_67_389 ();
 fill_1 FILLER_67_391 ();
 decap_12 FILLER_67_393 ();
 decap_12 FILLER_67_405 ();
 decap_12 FILLER_67_417 ();
 decap_12 FILLER_67_429 ();
 fill_4 FILLER_67_441 ();
 fill_2 FILLER_67_445 ();
 fill_1 FILLER_67_447 ();
 decap_12 FILLER_67_449 ();
 decap_12 FILLER_67_461 ();
 decap_12 FILLER_67_473 ();
 decap_12 FILLER_67_485 ();
 fill_4 FILLER_67_497 ();
 fill_2 FILLER_67_501 ();
 fill_1 FILLER_67_503 ();
 decap_12 FILLER_67_505 ();
 decap_12 FILLER_67_517 ();
 decap_12 FILLER_67_529 ();
 decap_12 FILLER_67_541 ();
 fill_4 FILLER_67_553 ();
 fill_2 FILLER_67_557 ();
 fill_1 FILLER_67_559 ();
 decap_12 FILLER_67_561 ();
 decap_12 FILLER_67_573 ();
 decap_12 FILLER_67_585 ();
 decap_12 FILLER_67_597 ();
 fill_4 FILLER_67_609 ();
 fill_2 FILLER_67_613 ();
 fill_1 FILLER_67_615 ();
 fill_8 FILLER_67_617 ();
 decap_12 FILLER_68_3 ();
 decap_12 FILLER_68_15 ();
 fill_1 FILLER_68_27 ();
 decap_12 FILLER_68_29 ();
 decap_12 FILLER_68_41 ();
 decap_12 FILLER_68_53 ();
 decap_12 FILLER_68_65 ();
 fill_4 FILLER_68_77 ();
 fill_2 FILLER_68_81 ();
 fill_1 FILLER_68_83 ();
 decap_12 FILLER_68_85 ();
 decap_12 FILLER_68_97 ();
 decap_12 FILLER_68_109 ();
 decap_12 FILLER_68_121 ();
 fill_4 FILLER_68_133 ();
 fill_2 FILLER_68_137 ();
 fill_1 FILLER_68_139 ();
 decap_12 FILLER_68_141 ();
 decap_12 FILLER_68_153 ();
 decap_12 FILLER_68_165 ();
 decap_12 FILLER_68_177 ();
 fill_4 FILLER_68_189 ();
 fill_2 FILLER_68_193 ();
 fill_1 FILLER_68_195 ();
 decap_12 FILLER_68_197 ();
 decap_12 FILLER_68_209 ();
 decap_12 FILLER_68_221 ();
 decap_12 FILLER_68_233 ();
 fill_4 FILLER_68_245 ();
 fill_2 FILLER_68_249 ();
 fill_1 FILLER_68_251 ();
 decap_12 FILLER_68_253 ();
 decap_12 FILLER_68_265 ();
 decap_12 FILLER_68_277 ();
 decap_12 FILLER_68_289 ();
 fill_4 FILLER_68_301 ();
 fill_2 FILLER_68_305 ();
 fill_1 FILLER_68_307 ();
 decap_12 FILLER_68_309 ();
 decap_12 FILLER_68_321 ();
 decap_12 FILLER_68_333 ();
 decap_12 FILLER_68_345 ();
 fill_4 FILLER_68_357 ();
 fill_2 FILLER_68_361 ();
 fill_1 FILLER_68_363 ();
 decap_12 FILLER_68_365 ();
 decap_12 FILLER_68_377 ();
 decap_12 FILLER_68_389 ();
 decap_12 FILLER_68_401 ();
 fill_4 FILLER_68_413 ();
 fill_2 FILLER_68_417 ();
 fill_1 FILLER_68_419 ();
 decap_12 FILLER_68_421 ();
 decap_12 FILLER_68_433 ();
 decap_12 FILLER_68_445 ();
 decap_12 FILLER_68_457 ();
 fill_4 FILLER_68_469 ();
 fill_2 FILLER_68_473 ();
 fill_1 FILLER_68_475 ();
 decap_12 FILLER_68_477 ();
 decap_12 FILLER_68_489 ();
 decap_12 FILLER_68_501 ();
 decap_12 FILLER_68_513 ();
 fill_4 FILLER_68_525 ();
 fill_2 FILLER_68_529 ();
 fill_1 FILLER_68_531 ();
 decap_12 FILLER_68_533 ();
 decap_12 FILLER_68_545 ();
 decap_12 FILLER_68_557 ();
 decap_12 FILLER_68_569 ();
 fill_4 FILLER_68_581 ();
 fill_2 FILLER_68_585 ();
 fill_1 FILLER_68_587 ();
 decap_12 FILLER_68_589 ();
 decap_12 FILLER_68_601 ();
 decap_12 FILLER_68_613 ();
 decap_12 FILLER_69_3 ();
 decap_12 FILLER_69_15 ();
 decap_12 FILLER_69_27 ();
 decap_12 FILLER_69_39 ();
 fill_4 FILLER_69_51 ();
 fill_1 FILLER_69_55 ();
 decap_12 FILLER_69_57 ();
 decap_12 FILLER_69_69 ();
 decap_12 FILLER_69_81 ();
 decap_12 FILLER_69_93 ();
 fill_4 FILLER_69_105 ();
 fill_2 FILLER_69_109 ();
 fill_1 FILLER_69_111 ();
 decap_12 FILLER_69_113 ();
 decap_12 FILLER_69_125 ();
 decap_12 FILLER_69_137 ();
 decap_12 FILLER_69_149 ();
 fill_4 FILLER_69_161 ();
 fill_2 FILLER_69_165 ();
 fill_1 FILLER_69_167 ();
 decap_12 FILLER_69_169 ();
 decap_12 FILLER_69_181 ();
 decap_12 FILLER_69_193 ();
 decap_12 FILLER_69_205 ();
 fill_4 FILLER_69_217 ();
 fill_2 FILLER_69_221 ();
 fill_1 FILLER_69_223 ();
 decap_12 FILLER_69_225 ();
 decap_12 FILLER_69_237 ();
 decap_12 FILLER_69_249 ();
 decap_12 FILLER_69_261 ();
 fill_4 FILLER_69_273 ();
 fill_2 FILLER_69_277 ();
 fill_1 FILLER_69_279 ();
 decap_12 FILLER_69_281 ();
 decap_12 FILLER_69_293 ();
 decap_12 FILLER_69_305 ();
 decap_12 FILLER_69_317 ();
 fill_4 FILLER_69_329 ();
 fill_2 FILLER_69_333 ();
 fill_1 FILLER_69_335 ();
 decap_12 FILLER_69_337 ();
 decap_12 FILLER_69_349 ();
 decap_12 FILLER_69_361 ();
 decap_12 FILLER_69_373 ();
 fill_4 FILLER_69_385 ();
 fill_2 FILLER_69_389 ();
 fill_1 FILLER_69_391 ();
 decap_12 FILLER_69_393 ();
 decap_12 FILLER_69_405 ();
 decap_12 FILLER_69_417 ();
 decap_12 FILLER_69_429 ();
 fill_4 FILLER_69_441 ();
 fill_2 FILLER_69_445 ();
 fill_1 FILLER_69_447 ();
 decap_12 FILLER_69_449 ();
 decap_12 FILLER_69_461 ();
 decap_12 FILLER_69_473 ();
 decap_12 FILLER_69_485 ();
 fill_4 FILLER_69_497 ();
 fill_2 FILLER_69_501 ();
 fill_1 FILLER_69_503 ();
 decap_12 FILLER_69_505 ();
 decap_12 FILLER_69_517 ();
 decap_12 FILLER_69_529 ();
 decap_12 FILLER_69_541 ();
 fill_4 FILLER_69_553 ();
 fill_2 FILLER_69_557 ();
 fill_1 FILLER_69_559 ();
 decap_12 FILLER_69_561 ();
 decap_12 FILLER_69_573 ();
 decap_12 FILLER_69_585 ();
 decap_12 FILLER_69_597 ();
 fill_4 FILLER_69_609 ();
 fill_2 FILLER_69_613 ();
 fill_1 FILLER_69_615 ();
 fill_8 FILLER_69_617 ();
 decap_12 FILLER_70_3 ();
 decap_12 FILLER_70_15 ();
 fill_1 FILLER_70_27 ();
 decap_12 FILLER_70_29 ();
 decap_12 FILLER_70_41 ();
 decap_12 FILLER_70_53 ();
 decap_12 FILLER_70_65 ();
 fill_4 FILLER_70_77 ();
 fill_2 FILLER_70_81 ();
 fill_1 FILLER_70_83 ();
 decap_12 FILLER_70_85 ();
 decap_12 FILLER_70_97 ();
 decap_12 FILLER_70_109 ();
 decap_12 FILLER_70_121 ();
 fill_4 FILLER_70_133 ();
 fill_2 FILLER_70_137 ();
 fill_1 FILLER_70_139 ();
 decap_12 FILLER_70_141 ();
 decap_12 FILLER_70_153 ();
 decap_12 FILLER_70_165 ();
 decap_12 FILLER_70_177 ();
 fill_4 FILLER_70_189 ();
 fill_2 FILLER_70_193 ();
 fill_1 FILLER_70_195 ();
 decap_12 FILLER_70_197 ();
 decap_12 FILLER_70_209 ();
 decap_12 FILLER_70_221 ();
 decap_12 FILLER_70_233 ();
 fill_4 FILLER_70_245 ();
 fill_2 FILLER_70_249 ();
 fill_1 FILLER_70_251 ();
 decap_12 FILLER_70_253 ();
 decap_12 FILLER_70_265 ();
 decap_12 FILLER_70_277 ();
 decap_12 FILLER_70_289 ();
 fill_4 FILLER_70_301 ();
 fill_2 FILLER_70_305 ();
 fill_1 FILLER_70_307 ();
 decap_12 FILLER_70_309 ();
 decap_12 FILLER_70_321 ();
 decap_12 FILLER_70_333 ();
 decap_12 FILLER_70_345 ();
 fill_4 FILLER_70_357 ();
 fill_2 FILLER_70_361 ();
 fill_1 FILLER_70_363 ();
 decap_12 FILLER_70_365 ();
 decap_12 FILLER_70_377 ();
 decap_12 FILLER_70_389 ();
 decap_12 FILLER_70_401 ();
 fill_4 FILLER_70_413 ();
 fill_2 FILLER_70_417 ();
 fill_1 FILLER_70_419 ();
 decap_12 FILLER_70_421 ();
 decap_12 FILLER_70_433 ();
 decap_12 FILLER_70_445 ();
 decap_12 FILLER_70_457 ();
 fill_4 FILLER_70_469 ();
 fill_2 FILLER_70_473 ();
 fill_1 FILLER_70_475 ();
 decap_12 FILLER_70_477 ();
 decap_12 FILLER_70_489 ();
 decap_12 FILLER_70_501 ();
 decap_12 FILLER_70_513 ();
 fill_4 FILLER_70_525 ();
 fill_2 FILLER_70_529 ();
 fill_1 FILLER_70_531 ();
 decap_12 FILLER_70_533 ();
 decap_12 FILLER_70_545 ();
 decap_12 FILLER_70_557 ();
 decap_12 FILLER_70_569 ();
 fill_4 FILLER_70_581 ();
 fill_2 FILLER_70_585 ();
 fill_1 FILLER_70_587 ();
 decap_12 FILLER_70_589 ();
 decap_12 FILLER_70_601 ();
 decap_12 FILLER_70_613 ();
 decap_12 FILLER_71_3 ();
 decap_12 FILLER_71_15 ();
 decap_12 FILLER_71_27 ();
 decap_12 FILLER_71_39 ();
 fill_4 FILLER_71_51 ();
 fill_1 FILLER_71_55 ();
 decap_12 FILLER_71_57 ();
 decap_12 FILLER_71_69 ();
 decap_12 FILLER_71_81 ();
 decap_12 FILLER_71_93 ();
 fill_4 FILLER_71_105 ();
 fill_2 FILLER_71_109 ();
 fill_1 FILLER_71_111 ();
 decap_12 FILLER_71_113 ();
 decap_12 FILLER_71_125 ();
 decap_12 FILLER_71_137 ();
 decap_12 FILLER_71_149 ();
 fill_4 FILLER_71_161 ();
 fill_2 FILLER_71_165 ();
 fill_1 FILLER_71_167 ();
 decap_12 FILLER_71_169 ();
 decap_12 FILLER_71_181 ();
 decap_12 FILLER_71_193 ();
 decap_12 FILLER_71_205 ();
 fill_4 FILLER_71_217 ();
 fill_2 FILLER_71_221 ();
 fill_1 FILLER_71_223 ();
 decap_12 FILLER_71_225 ();
 decap_12 FILLER_71_237 ();
 decap_12 FILLER_71_249 ();
 decap_12 FILLER_71_261 ();
 fill_4 FILLER_71_273 ();
 fill_2 FILLER_71_277 ();
 fill_1 FILLER_71_279 ();
 decap_12 FILLER_71_281 ();
 decap_12 FILLER_71_293 ();
 decap_12 FILLER_71_305 ();
 decap_12 FILLER_71_317 ();
 fill_4 FILLER_71_329 ();
 fill_2 FILLER_71_333 ();
 fill_1 FILLER_71_335 ();
 decap_12 FILLER_71_337 ();
 decap_12 FILLER_71_349 ();
 decap_12 FILLER_71_361 ();
 decap_12 FILLER_71_373 ();
 fill_4 FILLER_71_385 ();
 fill_2 FILLER_71_389 ();
 fill_1 FILLER_71_391 ();
 decap_12 FILLER_71_393 ();
 decap_12 FILLER_71_405 ();
 decap_12 FILLER_71_417 ();
 decap_12 FILLER_71_429 ();
 fill_4 FILLER_71_441 ();
 fill_2 FILLER_71_445 ();
 fill_1 FILLER_71_447 ();
 decap_12 FILLER_71_449 ();
 decap_12 FILLER_71_461 ();
 decap_12 FILLER_71_473 ();
 decap_12 FILLER_71_485 ();
 fill_4 FILLER_71_497 ();
 fill_2 FILLER_71_501 ();
 fill_1 FILLER_71_503 ();
 decap_12 FILLER_71_505 ();
 decap_12 FILLER_71_517 ();
 decap_12 FILLER_71_529 ();
 decap_12 FILLER_71_541 ();
 fill_4 FILLER_71_553 ();
 fill_2 FILLER_71_557 ();
 fill_1 FILLER_71_559 ();
 decap_12 FILLER_71_561 ();
 decap_12 FILLER_71_573 ();
 decap_12 FILLER_71_585 ();
 decap_12 FILLER_71_597 ();
 fill_4 FILLER_71_609 ();
 fill_2 FILLER_71_613 ();
 fill_1 FILLER_71_615 ();
 fill_8 FILLER_71_617 ();
 decap_12 FILLER_72_3 ();
 decap_12 FILLER_72_15 ();
 fill_1 FILLER_72_27 ();
 decap_12 FILLER_72_29 ();
 decap_12 FILLER_72_41 ();
 decap_12 FILLER_72_53 ();
 decap_12 FILLER_72_65 ();
 fill_4 FILLER_72_77 ();
 fill_2 FILLER_72_81 ();
 fill_1 FILLER_72_83 ();
 decap_12 FILLER_72_85 ();
 decap_12 FILLER_72_97 ();
 decap_12 FILLER_72_109 ();
 decap_12 FILLER_72_121 ();
 fill_4 FILLER_72_133 ();
 fill_2 FILLER_72_137 ();
 fill_1 FILLER_72_139 ();
 decap_12 FILLER_72_141 ();
 decap_12 FILLER_72_153 ();
 decap_12 FILLER_72_165 ();
 decap_12 FILLER_72_177 ();
 fill_4 FILLER_72_189 ();
 fill_2 FILLER_72_193 ();
 fill_1 FILLER_72_195 ();
 decap_12 FILLER_72_197 ();
 decap_12 FILLER_72_209 ();
 decap_12 FILLER_72_221 ();
 decap_12 FILLER_72_233 ();
 fill_4 FILLER_72_245 ();
 fill_2 FILLER_72_249 ();
 fill_1 FILLER_72_251 ();
 decap_12 FILLER_72_253 ();
 decap_12 FILLER_72_265 ();
 decap_12 FILLER_72_277 ();
 decap_12 FILLER_72_289 ();
 fill_4 FILLER_72_301 ();
 fill_2 FILLER_72_305 ();
 fill_1 FILLER_72_307 ();
 decap_12 FILLER_72_309 ();
 decap_12 FILLER_72_321 ();
 decap_12 FILLER_72_333 ();
 decap_12 FILLER_72_345 ();
 fill_4 FILLER_72_357 ();
 fill_2 FILLER_72_361 ();
 fill_1 FILLER_72_363 ();
 decap_12 FILLER_72_365 ();
 decap_12 FILLER_72_377 ();
 decap_12 FILLER_72_389 ();
 decap_12 FILLER_72_401 ();
 fill_4 FILLER_72_413 ();
 fill_2 FILLER_72_417 ();
 fill_1 FILLER_72_419 ();
 decap_12 FILLER_72_421 ();
 decap_12 FILLER_72_433 ();
 decap_12 FILLER_72_445 ();
 decap_12 FILLER_72_457 ();
 fill_4 FILLER_72_469 ();
 fill_2 FILLER_72_473 ();
 fill_1 FILLER_72_475 ();
 decap_12 FILLER_72_477 ();
 decap_12 FILLER_72_489 ();
 decap_12 FILLER_72_501 ();
 decap_12 FILLER_72_513 ();
 fill_4 FILLER_72_525 ();
 fill_2 FILLER_72_529 ();
 fill_1 FILLER_72_531 ();
 decap_12 FILLER_72_533 ();
 decap_12 FILLER_72_545 ();
 decap_12 FILLER_72_557 ();
 decap_12 FILLER_72_569 ();
 fill_4 FILLER_72_581 ();
 fill_2 FILLER_72_585 ();
 fill_1 FILLER_72_587 ();
 decap_12 FILLER_72_589 ();
 decap_12 FILLER_72_601 ();
 decap_12 FILLER_72_613 ();
 decap_12 FILLER_73_3 ();
 decap_12 FILLER_73_15 ();
 decap_12 FILLER_73_27 ();
 decap_12 FILLER_73_39 ();
 fill_4 FILLER_73_51 ();
 fill_1 FILLER_73_55 ();
 decap_12 FILLER_73_57 ();
 decap_12 FILLER_73_69 ();
 decap_12 FILLER_73_81 ();
 decap_12 FILLER_73_93 ();
 fill_4 FILLER_73_105 ();
 fill_2 FILLER_73_109 ();
 fill_1 FILLER_73_111 ();
 decap_12 FILLER_73_113 ();
 decap_12 FILLER_73_125 ();
 decap_12 FILLER_73_137 ();
 decap_12 FILLER_73_149 ();
 fill_4 FILLER_73_161 ();
 fill_2 FILLER_73_165 ();
 fill_1 FILLER_73_167 ();
 decap_12 FILLER_73_169 ();
 decap_12 FILLER_73_181 ();
 decap_12 FILLER_73_193 ();
 decap_12 FILLER_73_205 ();
 fill_4 FILLER_73_217 ();
 fill_2 FILLER_73_221 ();
 fill_1 FILLER_73_223 ();
 decap_12 FILLER_73_225 ();
 decap_12 FILLER_73_237 ();
 decap_12 FILLER_73_249 ();
 decap_12 FILLER_73_261 ();
 fill_4 FILLER_73_273 ();
 fill_2 FILLER_73_277 ();
 fill_1 FILLER_73_279 ();
 decap_12 FILLER_73_281 ();
 decap_12 FILLER_73_293 ();
 decap_12 FILLER_73_305 ();
 decap_12 FILLER_73_317 ();
 fill_4 FILLER_73_329 ();
 fill_2 FILLER_73_333 ();
 fill_1 FILLER_73_335 ();
 decap_12 FILLER_73_337 ();
 decap_12 FILLER_73_349 ();
 decap_12 FILLER_73_361 ();
 decap_12 FILLER_73_373 ();
 fill_4 FILLER_73_385 ();
 fill_2 FILLER_73_389 ();
 fill_1 FILLER_73_391 ();
 decap_12 FILLER_73_393 ();
 decap_12 FILLER_73_405 ();
 decap_12 FILLER_73_417 ();
 decap_12 FILLER_73_429 ();
 fill_4 FILLER_73_441 ();
 fill_2 FILLER_73_445 ();
 fill_1 FILLER_73_447 ();
 decap_12 FILLER_73_449 ();
 decap_12 FILLER_73_461 ();
 decap_12 FILLER_73_473 ();
 decap_12 FILLER_73_485 ();
 fill_4 FILLER_73_497 ();
 fill_2 FILLER_73_501 ();
 fill_1 FILLER_73_503 ();
 decap_12 FILLER_73_505 ();
 decap_12 FILLER_73_517 ();
 decap_12 FILLER_73_529 ();
 decap_12 FILLER_73_541 ();
 fill_4 FILLER_73_553 ();
 fill_2 FILLER_73_557 ();
 fill_1 FILLER_73_559 ();
 decap_12 FILLER_73_561 ();
 decap_12 FILLER_73_573 ();
 decap_12 FILLER_73_585 ();
 decap_12 FILLER_73_597 ();
 fill_4 FILLER_73_609 ();
 fill_2 FILLER_73_613 ();
 fill_1 FILLER_73_615 ();
 fill_8 FILLER_73_617 ();
 decap_12 FILLER_74_3 ();
 decap_12 FILLER_74_15 ();
 fill_1 FILLER_74_27 ();
 decap_12 FILLER_74_29 ();
 decap_12 FILLER_74_41 ();
 decap_12 FILLER_74_53 ();
 decap_12 FILLER_74_65 ();
 fill_4 FILLER_74_77 ();
 fill_2 FILLER_74_81 ();
 fill_1 FILLER_74_83 ();
 decap_12 FILLER_74_85 ();
 decap_12 FILLER_74_97 ();
 decap_12 FILLER_74_109 ();
 decap_12 FILLER_74_121 ();
 fill_4 FILLER_74_133 ();
 fill_2 FILLER_74_137 ();
 fill_1 FILLER_74_139 ();
 decap_12 FILLER_74_141 ();
 decap_12 FILLER_74_153 ();
 decap_12 FILLER_74_165 ();
 decap_12 FILLER_74_177 ();
 fill_4 FILLER_74_189 ();
 fill_2 FILLER_74_193 ();
 fill_1 FILLER_74_195 ();
 decap_12 FILLER_74_197 ();
 decap_12 FILLER_74_209 ();
 decap_12 FILLER_74_221 ();
 decap_12 FILLER_74_233 ();
 fill_4 FILLER_74_245 ();
 fill_2 FILLER_74_249 ();
 fill_1 FILLER_74_251 ();
 decap_12 FILLER_74_253 ();
 decap_12 FILLER_74_265 ();
 decap_12 FILLER_74_277 ();
 decap_12 FILLER_74_289 ();
 fill_4 FILLER_74_301 ();
 fill_2 FILLER_74_305 ();
 fill_1 FILLER_74_307 ();
 decap_12 FILLER_74_309 ();
 decap_12 FILLER_74_321 ();
 decap_12 FILLER_74_333 ();
 decap_12 FILLER_74_345 ();
 fill_4 FILLER_74_357 ();
 fill_2 FILLER_74_361 ();
 fill_1 FILLER_74_363 ();
 decap_12 FILLER_74_365 ();
 decap_12 FILLER_74_377 ();
 decap_12 FILLER_74_389 ();
 decap_12 FILLER_74_401 ();
 fill_4 FILLER_74_413 ();
 fill_2 FILLER_74_417 ();
 fill_1 FILLER_74_419 ();
 decap_12 FILLER_74_421 ();
 decap_12 FILLER_74_433 ();
 decap_12 FILLER_74_445 ();
 decap_12 FILLER_74_457 ();
 fill_4 FILLER_74_469 ();
 fill_2 FILLER_74_473 ();
 fill_1 FILLER_74_475 ();
 decap_12 FILLER_74_477 ();
 decap_12 FILLER_74_489 ();
 decap_12 FILLER_74_501 ();
 decap_12 FILLER_74_513 ();
 fill_4 FILLER_74_525 ();
 fill_2 FILLER_74_529 ();
 fill_1 FILLER_74_531 ();
 decap_12 FILLER_74_533 ();
 decap_12 FILLER_74_545 ();
 decap_12 FILLER_74_557 ();
 decap_12 FILLER_74_569 ();
 fill_4 FILLER_74_581 ();
 fill_2 FILLER_74_585 ();
 fill_1 FILLER_74_587 ();
 decap_12 FILLER_74_589 ();
 decap_12 FILLER_74_601 ();
 decap_12 FILLER_74_613 ();
 decap_12 FILLER_75_3 ();
 decap_12 FILLER_75_15 ();
 decap_12 FILLER_75_27 ();
 decap_12 FILLER_75_39 ();
 fill_4 FILLER_75_51 ();
 fill_1 FILLER_75_55 ();
 decap_12 FILLER_75_57 ();
 decap_12 FILLER_75_69 ();
 decap_12 FILLER_75_81 ();
 decap_12 FILLER_75_93 ();
 fill_4 FILLER_75_105 ();
 fill_2 FILLER_75_109 ();
 fill_1 FILLER_75_111 ();
 decap_12 FILLER_75_113 ();
 decap_12 FILLER_75_125 ();
 decap_12 FILLER_75_137 ();
 decap_12 FILLER_75_149 ();
 fill_4 FILLER_75_161 ();
 fill_2 FILLER_75_165 ();
 fill_1 FILLER_75_167 ();
 decap_12 FILLER_75_169 ();
 decap_12 FILLER_75_181 ();
 decap_12 FILLER_75_193 ();
 decap_12 FILLER_75_205 ();
 fill_4 FILLER_75_217 ();
 fill_2 FILLER_75_221 ();
 fill_1 FILLER_75_223 ();
 decap_12 FILLER_75_225 ();
 decap_12 FILLER_75_237 ();
 decap_12 FILLER_75_249 ();
 decap_12 FILLER_75_261 ();
 fill_4 FILLER_75_273 ();
 fill_2 FILLER_75_277 ();
 fill_1 FILLER_75_279 ();
 decap_12 FILLER_75_281 ();
 decap_12 FILLER_75_293 ();
 decap_12 FILLER_75_305 ();
 decap_12 FILLER_75_317 ();
 fill_4 FILLER_75_329 ();
 fill_2 FILLER_75_333 ();
 fill_1 FILLER_75_335 ();
 decap_12 FILLER_75_337 ();
 decap_12 FILLER_75_349 ();
 decap_12 FILLER_75_361 ();
 decap_12 FILLER_75_373 ();
 fill_4 FILLER_75_385 ();
 fill_2 FILLER_75_389 ();
 fill_1 FILLER_75_391 ();
 decap_12 FILLER_75_393 ();
 decap_12 FILLER_75_405 ();
 decap_12 FILLER_75_417 ();
 decap_12 FILLER_75_429 ();
 fill_4 FILLER_75_441 ();
 fill_2 FILLER_75_445 ();
 fill_1 FILLER_75_447 ();
 decap_12 FILLER_75_449 ();
 decap_12 FILLER_75_461 ();
 decap_12 FILLER_75_473 ();
 decap_12 FILLER_75_485 ();
 fill_4 FILLER_75_497 ();
 fill_2 FILLER_75_501 ();
 fill_1 FILLER_75_503 ();
 decap_12 FILLER_75_505 ();
 decap_12 FILLER_75_517 ();
 decap_12 FILLER_75_529 ();
 decap_12 FILLER_75_541 ();
 fill_4 FILLER_75_553 ();
 fill_2 FILLER_75_557 ();
 fill_1 FILLER_75_559 ();
 decap_12 FILLER_75_561 ();
 decap_12 FILLER_75_573 ();
 decap_12 FILLER_75_585 ();
 decap_12 FILLER_75_597 ();
 fill_4 FILLER_75_609 ();
 fill_2 FILLER_75_613 ();
 fill_1 FILLER_75_615 ();
 fill_8 FILLER_75_617 ();
 decap_12 FILLER_76_3 ();
 decap_12 FILLER_76_15 ();
 fill_1 FILLER_76_27 ();
 decap_12 FILLER_76_29 ();
 decap_12 FILLER_76_41 ();
 decap_12 FILLER_76_53 ();
 decap_12 FILLER_76_65 ();
 fill_4 FILLER_76_77 ();
 fill_2 FILLER_76_81 ();
 fill_1 FILLER_76_83 ();
 decap_12 FILLER_76_85 ();
 decap_12 FILLER_76_97 ();
 decap_12 FILLER_76_109 ();
 decap_12 FILLER_76_121 ();
 fill_4 FILLER_76_133 ();
 fill_2 FILLER_76_137 ();
 fill_1 FILLER_76_139 ();
 decap_12 FILLER_76_141 ();
 decap_12 FILLER_76_153 ();
 decap_12 FILLER_76_165 ();
 decap_12 FILLER_76_177 ();
 fill_4 FILLER_76_189 ();
 fill_2 FILLER_76_193 ();
 fill_1 FILLER_76_195 ();
 decap_12 FILLER_76_197 ();
 decap_12 FILLER_76_209 ();
 decap_12 FILLER_76_221 ();
 decap_12 FILLER_76_233 ();
 fill_4 FILLER_76_245 ();
 fill_2 FILLER_76_249 ();
 fill_1 FILLER_76_251 ();
 decap_12 FILLER_76_253 ();
 decap_12 FILLER_76_265 ();
 decap_12 FILLER_76_277 ();
 decap_12 FILLER_76_289 ();
 fill_4 FILLER_76_301 ();
 fill_2 FILLER_76_305 ();
 fill_1 FILLER_76_307 ();
 decap_12 FILLER_76_309 ();
 decap_12 FILLER_76_321 ();
 decap_12 FILLER_76_333 ();
 decap_12 FILLER_76_345 ();
 fill_4 FILLER_76_357 ();
 fill_2 FILLER_76_361 ();
 fill_1 FILLER_76_363 ();
 decap_12 FILLER_76_365 ();
 decap_12 FILLER_76_377 ();
 decap_12 FILLER_76_389 ();
 decap_12 FILLER_76_401 ();
 fill_4 FILLER_76_413 ();
 fill_2 FILLER_76_417 ();
 fill_1 FILLER_76_419 ();
 decap_12 FILLER_76_421 ();
 decap_12 FILLER_76_433 ();
 decap_12 FILLER_76_445 ();
 decap_12 FILLER_76_457 ();
 fill_4 FILLER_76_469 ();
 fill_2 FILLER_76_473 ();
 fill_1 FILLER_76_475 ();
 decap_12 FILLER_76_477 ();
 decap_12 FILLER_76_489 ();
 decap_12 FILLER_76_501 ();
 decap_12 FILLER_76_513 ();
 fill_4 FILLER_76_525 ();
 fill_2 FILLER_76_529 ();
 fill_1 FILLER_76_531 ();
 decap_12 FILLER_76_533 ();
 decap_12 FILLER_76_545 ();
 decap_12 FILLER_76_557 ();
 decap_12 FILLER_76_569 ();
 fill_4 FILLER_76_581 ();
 fill_2 FILLER_76_585 ();
 fill_1 FILLER_76_587 ();
 decap_12 FILLER_76_589 ();
 decap_12 FILLER_76_601 ();
 decap_12 FILLER_76_613 ();
 decap_12 FILLER_77_3 ();
 decap_12 FILLER_77_15 ();
 decap_12 FILLER_77_27 ();
 decap_12 FILLER_77_39 ();
 fill_4 FILLER_77_51 ();
 fill_1 FILLER_77_55 ();
 decap_12 FILLER_77_57 ();
 decap_12 FILLER_77_69 ();
 decap_12 FILLER_77_81 ();
 decap_12 FILLER_77_93 ();
 fill_4 FILLER_77_105 ();
 fill_2 FILLER_77_109 ();
 fill_1 FILLER_77_111 ();
 decap_12 FILLER_77_113 ();
 decap_12 FILLER_77_125 ();
 decap_12 FILLER_77_137 ();
 decap_12 FILLER_77_149 ();
 fill_4 FILLER_77_161 ();
 fill_2 FILLER_77_165 ();
 fill_1 FILLER_77_167 ();
 decap_12 FILLER_77_169 ();
 decap_12 FILLER_77_181 ();
 decap_12 FILLER_77_193 ();
 decap_12 FILLER_77_205 ();
 fill_4 FILLER_77_217 ();
 fill_2 FILLER_77_221 ();
 fill_1 FILLER_77_223 ();
 decap_12 FILLER_77_225 ();
 decap_12 FILLER_77_237 ();
 decap_12 FILLER_77_249 ();
 decap_12 FILLER_77_261 ();
 fill_4 FILLER_77_273 ();
 fill_2 FILLER_77_277 ();
 fill_1 FILLER_77_279 ();
 decap_12 FILLER_77_281 ();
 decap_12 FILLER_77_293 ();
 decap_12 FILLER_77_305 ();
 decap_12 FILLER_77_317 ();
 fill_4 FILLER_77_329 ();
 fill_2 FILLER_77_333 ();
 fill_1 FILLER_77_335 ();
 decap_12 FILLER_77_337 ();
 decap_12 FILLER_77_349 ();
 decap_12 FILLER_77_361 ();
 decap_12 FILLER_77_373 ();
 fill_4 FILLER_77_385 ();
 fill_2 FILLER_77_389 ();
 fill_1 FILLER_77_391 ();
 decap_12 FILLER_77_393 ();
 decap_12 FILLER_77_405 ();
 decap_12 FILLER_77_417 ();
 decap_12 FILLER_77_429 ();
 fill_4 FILLER_77_441 ();
 fill_2 FILLER_77_445 ();
 fill_1 FILLER_77_447 ();
 decap_12 FILLER_77_449 ();
 decap_12 FILLER_77_461 ();
 decap_12 FILLER_77_473 ();
 decap_12 FILLER_77_485 ();
 fill_4 FILLER_77_497 ();
 fill_2 FILLER_77_501 ();
 fill_1 FILLER_77_503 ();
 decap_12 FILLER_77_505 ();
 decap_12 FILLER_77_517 ();
 decap_12 FILLER_77_529 ();
 decap_12 FILLER_77_541 ();
 fill_4 FILLER_77_553 ();
 fill_2 FILLER_77_557 ();
 fill_1 FILLER_77_559 ();
 decap_12 FILLER_77_561 ();
 decap_12 FILLER_77_573 ();
 decap_12 FILLER_77_585 ();
 decap_12 FILLER_77_597 ();
 fill_4 FILLER_77_609 ();
 fill_2 FILLER_77_613 ();
 fill_1 FILLER_77_615 ();
 fill_8 FILLER_77_617 ();
 decap_12 FILLER_78_3 ();
 decap_12 FILLER_78_15 ();
 fill_1 FILLER_78_27 ();
 decap_12 FILLER_78_29 ();
 decap_12 FILLER_78_41 ();
 decap_12 FILLER_78_53 ();
 decap_12 FILLER_78_65 ();
 fill_4 FILLER_78_77 ();
 fill_2 FILLER_78_81 ();
 fill_1 FILLER_78_83 ();
 decap_12 FILLER_78_85 ();
 decap_12 FILLER_78_97 ();
 decap_12 FILLER_78_109 ();
 decap_12 FILLER_78_121 ();
 fill_4 FILLER_78_133 ();
 fill_2 FILLER_78_137 ();
 fill_1 FILLER_78_139 ();
 decap_12 FILLER_78_141 ();
 decap_12 FILLER_78_153 ();
 decap_12 FILLER_78_165 ();
 decap_12 FILLER_78_177 ();
 fill_4 FILLER_78_189 ();
 fill_2 FILLER_78_193 ();
 fill_1 FILLER_78_195 ();
 decap_12 FILLER_78_197 ();
 decap_12 FILLER_78_209 ();
 decap_12 FILLER_78_221 ();
 decap_12 FILLER_78_233 ();
 fill_4 FILLER_78_245 ();
 fill_2 FILLER_78_249 ();
 fill_1 FILLER_78_251 ();
 decap_12 FILLER_78_253 ();
 decap_12 FILLER_78_265 ();
 decap_12 FILLER_78_277 ();
 decap_12 FILLER_78_289 ();
 fill_4 FILLER_78_301 ();
 fill_2 FILLER_78_305 ();
 fill_1 FILLER_78_307 ();
 decap_12 FILLER_78_309 ();
 decap_12 FILLER_78_321 ();
 decap_12 FILLER_78_333 ();
 decap_12 FILLER_78_345 ();
 fill_4 FILLER_78_357 ();
 fill_2 FILLER_78_361 ();
 fill_1 FILLER_78_363 ();
 decap_12 FILLER_78_365 ();
 decap_12 FILLER_78_377 ();
 decap_12 FILLER_78_389 ();
 decap_12 FILLER_78_401 ();
 fill_4 FILLER_78_413 ();
 fill_2 FILLER_78_417 ();
 fill_1 FILLER_78_419 ();
 decap_12 FILLER_78_421 ();
 decap_12 FILLER_78_433 ();
 decap_12 FILLER_78_445 ();
 decap_12 FILLER_78_457 ();
 fill_4 FILLER_78_469 ();
 fill_2 FILLER_78_473 ();
 fill_1 FILLER_78_475 ();
 decap_12 FILLER_78_477 ();
 decap_12 FILLER_78_489 ();
 decap_12 FILLER_78_501 ();
 decap_12 FILLER_78_513 ();
 fill_4 FILLER_78_525 ();
 fill_2 FILLER_78_529 ();
 fill_1 FILLER_78_531 ();
 decap_12 FILLER_78_533 ();
 decap_12 FILLER_78_545 ();
 decap_12 FILLER_78_557 ();
 decap_12 FILLER_78_569 ();
 fill_4 FILLER_78_581 ();
 fill_2 FILLER_78_585 ();
 fill_1 FILLER_78_587 ();
 decap_12 FILLER_78_589 ();
 decap_12 FILLER_78_601 ();
 decap_12 FILLER_78_613 ();
 decap_12 FILLER_79_3 ();
 decap_12 FILLER_79_15 ();
 decap_12 FILLER_79_27 ();
 decap_12 FILLER_79_39 ();
 fill_4 FILLER_79_51 ();
 fill_1 FILLER_79_55 ();
 decap_12 FILLER_79_57 ();
 decap_12 FILLER_79_69 ();
 decap_12 FILLER_79_81 ();
 decap_12 FILLER_79_93 ();
 fill_4 FILLER_79_105 ();
 fill_2 FILLER_79_109 ();
 fill_1 FILLER_79_111 ();
 decap_12 FILLER_79_113 ();
 decap_12 FILLER_79_125 ();
 decap_12 FILLER_79_137 ();
 decap_12 FILLER_79_149 ();
 fill_4 FILLER_79_161 ();
 fill_2 FILLER_79_165 ();
 fill_1 FILLER_79_167 ();
 decap_12 FILLER_79_169 ();
 decap_12 FILLER_79_181 ();
 decap_12 FILLER_79_193 ();
 decap_12 FILLER_79_205 ();
 fill_4 FILLER_79_217 ();
 fill_2 FILLER_79_221 ();
 fill_1 FILLER_79_223 ();
 decap_12 FILLER_79_225 ();
 decap_12 FILLER_79_237 ();
 decap_12 FILLER_79_249 ();
 decap_12 FILLER_79_261 ();
 fill_4 FILLER_79_273 ();
 fill_2 FILLER_79_277 ();
 fill_1 FILLER_79_279 ();
 decap_12 FILLER_79_281 ();
 decap_12 FILLER_79_293 ();
 decap_12 FILLER_79_305 ();
 decap_12 FILLER_79_317 ();
 fill_4 FILLER_79_329 ();
 fill_2 FILLER_79_333 ();
 fill_1 FILLER_79_335 ();
 decap_12 FILLER_79_337 ();
 decap_12 FILLER_79_349 ();
 decap_12 FILLER_79_361 ();
 decap_12 FILLER_79_373 ();
 fill_4 FILLER_79_385 ();
 fill_2 FILLER_79_389 ();
 fill_1 FILLER_79_391 ();
 decap_12 FILLER_79_393 ();
 decap_12 FILLER_79_405 ();
 decap_12 FILLER_79_417 ();
 decap_12 FILLER_79_429 ();
 fill_4 FILLER_79_441 ();
 fill_2 FILLER_79_445 ();
 fill_1 FILLER_79_447 ();
 decap_12 FILLER_79_449 ();
 decap_12 FILLER_79_461 ();
 decap_12 FILLER_79_473 ();
 decap_12 FILLER_79_485 ();
 fill_4 FILLER_79_497 ();
 fill_2 FILLER_79_501 ();
 fill_1 FILLER_79_503 ();
 decap_12 FILLER_79_505 ();
 decap_12 FILLER_79_517 ();
 decap_12 FILLER_79_529 ();
 decap_12 FILLER_79_541 ();
 fill_4 FILLER_79_553 ();
 fill_2 FILLER_79_557 ();
 fill_1 FILLER_79_559 ();
 decap_12 FILLER_79_561 ();
 decap_12 FILLER_79_573 ();
 decap_12 FILLER_79_585 ();
 decap_12 FILLER_79_597 ();
 fill_4 FILLER_79_609 ();
 fill_2 FILLER_79_613 ();
 fill_1 FILLER_79_615 ();
 fill_8 FILLER_79_617 ();
 decap_12 FILLER_80_3 ();
 decap_12 FILLER_80_15 ();
 fill_1 FILLER_80_27 ();
 decap_12 FILLER_80_29 ();
 decap_12 FILLER_80_41 ();
 decap_12 FILLER_80_53 ();
 decap_12 FILLER_80_65 ();
 fill_4 FILLER_80_77 ();
 fill_2 FILLER_80_81 ();
 fill_1 FILLER_80_83 ();
 decap_12 FILLER_80_85 ();
 decap_12 FILLER_80_97 ();
 decap_12 FILLER_80_109 ();
 decap_12 FILLER_80_121 ();
 fill_4 FILLER_80_133 ();
 fill_2 FILLER_80_137 ();
 fill_1 FILLER_80_139 ();
 decap_12 FILLER_80_141 ();
 decap_12 FILLER_80_153 ();
 decap_12 FILLER_80_165 ();
 decap_12 FILLER_80_177 ();
 fill_4 FILLER_80_189 ();
 fill_2 FILLER_80_193 ();
 fill_1 FILLER_80_195 ();
 decap_12 FILLER_80_197 ();
 decap_12 FILLER_80_209 ();
 decap_12 FILLER_80_221 ();
 decap_12 FILLER_80_233 ();
 fill_4 FILLER_80_245 ();
 fill_2 FILLER_80_249 ();
 fill_1 FILLER_80_251 ();
 decap_12 FILLER_80_253 ();
 decap_12 FILLER_80_265 ();
 decap_12 FILLER_80_277 ();
 decap_12 FILLER_80_289 ();
 fill_4 FILLER_80_301 ();
 fill_2 FILLER_80_305 ();
 fill_1 FILLER_80_307 ();
 decap_12 FILLER_80_309 ();
 decap_12 FILLER_80_321 ();
 decap_12 FILLER_80_333 ();
 decap_12 FILLER_80_345 ();
 fill_4 FILLER_80_357 ();
 fill_2 FILLER_80_361 ();
 fill_1 FILLER_80_363 ();
 decap_12 FILLER_80_365 ();
 decap_12 FILLER_80_377 ();
 decap_12 FILLER_80_389 ();
 decap_12 FILLER_80_401 ();
 fill_4 FILLER_80_413 ();
 fill_2 FILLER_80_417 ();
 fill_1 FILLER_80_419 ();
 decap_12 FILLER_80_421 ();
 decap_12 FILLER_80_433 ();
 decap_12 FILLER_80_445 ();
 decap_12 FILLER_80_457 ();
 fill_4 FILLER_80_469 ();
 fill_2 FILLER_80_473 ();
 fill_1 FILLER_80_475 ();
 decap_12 FILLER_80_477 ();
 decap_12 FILLER_80_489 ();
 decap_12 FILLER_80_501 ();
 decap_12 FILLER_80_513 ();
 fill_4 FILLER_80_525 ();
 fill_2 FILLER_80_529 ();
 fill_1 FILLER_80_531 ();
 decap_12 FILLER_80_533 ();
 decap_12 FILLER_80_545 ();
 decap_12 FILLER_80_557 ();
 decap_12 FILLER_80_569 ();
 fill_4 FILLER_80_581 ();
 fill_2 FILLER_80_585 ();
 fill_1 FILLER_80_587 ();
 decap_12 FILLER_80_589 ();
 decap_12 FILLER_80_601 ();
 decap_12 FILLER_80_613 ();
 decap_12 FILLER_81_3 ();
 decap_12 FILLER_81_15 ();
 decap_12 FILLER_81_27 ();
 decap_12 FILLER_81_39 ();
 fill_4 FILLER_81_51 ();
 fill_1 FILLER_81_55 ();
 decap_12 FILLER_81_57 ();
 decap_12 FILLER_81_69 ();
 decap_12 FILLER_81_81 ();
 decap_12 FILLER_81_93 ();
 fill_4 FILLER_81_105 ();
 fill_2 FILLER_81_109 ();
 fill_1 FILLER_81_111 ();
 decap_12 FILLER_81_113 ();
 decap_12 FILLER_81_125 ();
 decap_12 FILLER_81_137 ();
 decap_12 FILLER_81_149 ();
 fill_4 FILLER_81_161 ();
 fill_2 FILLER_81_165 ();
 fill_1 FILLER_81_167 ();
 decap_12 FILLER_81_169 ();
 decap_12 FILLER_81_181 ();
 decap_12 FILLER_81_193 ();
 decap_12 FILLER_81_205 ();
 fill_4 FILLER_81_217 ();
 fill_2 FILLER_81_221 ();
 fill_1 FILLER_81_223 ();
 decap_12 FILLER_81_225 ();
 decap_12 FILLER_81_237 ();
 decap_12 FILLER_81_249 ();
 decap_12 FILLER_81_261 ();
 fill_4 FILLER_81_273 ();
 fill_2 FILLER_81_277 ();
 fill_1 FILLER_81_279 ();
 decap_12 FILLER_81_281 ();
 decap_12 FILLER_81_293 ();
 decap_12 FILLER_81_305 ();
 decap_12 FILLER_81_317 ();
 fill_4 FILLER_81_329 ();
 fill_2 FILLER_81_333 ();
 fill_1 FILLER_81_335 ();
 decap_12 FILLER_81_337 ();
 decap_12 FILLER_81_349 ();
 decap_12 FILLER_81_361 ();
 decap_12 FILLER_81_373 ();
 fill_4 FILLER_81_385 ();
 fill_2 FILLER_81_389 ();
 fill_1 FILLER_81_391 ();
 decap_12 FILLER_81_393 ();
 decap_12 FILLER_81_405 ();
 decap_12 FILLER_81_417 ();
 decap_12 FILLER_81_429 ();
 fill_4 FILLER_81_441 ();
 fill_2 FILLER_81_445 ();
 fill_1 FILLER_81_447 ();
 decap_12 FILLER_81_449 ();
 decap_12 FILLER_81_461 ();
 decap_12 FILLER_81_473 ();
 decap_12 FILLER_81_485 ();
 fill_4 FILLER_81_497 ();
 fill_2 FILLER_81_501 ();
 fill_1 FILLER_81_503 ();
 decap_12 FILLER_81_505 ();
 decap_12 FILLER_81_517 ();
 decap_12 FILLER_81_529 ();
 decap_12 FILLER_81_541 ();
 fill_4 FILLER_81_553 ();
 fill_2 FILLER_81_557 ();
 fill_1 FILLER_81_559 ();
 decap_12 FILLER_81_561 ();
 decap_12 FILLER_81_573 ();
 decap_12 FILLER_81_585 ();
 decap_12 FILLER_81_597 ();
 fill_4 FILLER_81_609 ();
 fill_2 FILLER_81_613 ();
 fill_1 FILLER_81_615 ();
 fill_8 FILLER_81_617 ();
 decap_12 FILLER_82_3 ();
 decap_12 FILLER_82_15 ();
 fill_1 FILLER_82_27 ();
 decap_12 FILLER_82_29 ();
 decap_12 FILLER_82_41 ();
 decap_12 FILLER_82_53 ();
 decap_12 FILLER_82_65 ();
 fill_4 FILLER_82_77 ();
 fill_2 FILLER_82_81 ();
 fill_1 FILLER_82_83 ();
 decap_12 FILLER_82_85 ();
 decap_12 FILLER_82_97 ();
 decap_12 FILLER_82_109 ();
 decap_12 FILLER_82_121 ();
 fill_4 FILLER_82_133 ();
 fill_2 FILLER_82_137 ();
 fill_1 FILLER_82_139 ();
 decap_12 FILLER_82_141 ();
 decap_12 FILLER_82_153 ();
 decap_12 FILLER_82_165 ();
 decap_12 FILLER_82_177 ();
 fill_4 FILLER_82_189 ();
 fill_2 FILLER_82_193 ();
 fill_1 FILLER_82_195 ();
 decap_12 FILLER_82_197 ();
 decap_12 FILLER_82_209 ();
 decap_12 FILLER_82_221 ();
 decap_12 FILLER_82_233 ();
 fill_4 FILLER_82_245 ();
 fill_2 FILLER_82_249 ();
 fill_1 FILLER_82_251 ();
 decap_12 FILLER_82_253 ();
 decap_12 FILLER_82_265 ();
 decap_12 FILLER_82_277 ();
 decap_12 FILLER_82_289 ();
 fill_4 FILLER_82_301 ();
 fill_2 FILLER_82_305 ();
 fill_1 FILLER_82_307 ();
 decap_12 FILLER_82_309 ();
 decap_12 FILLER_82_321 ();
 decap_12 FILLER_82_333 ();
 decap_12 FILLER_82_345 ();
 fill_4 FILLER_82_357 ();
 fill_2 FILLER_82_361 ();
 fill_1 FILLER_82_363 ();
 decap_12 FILLER_82_365 ();
 decap_12 FILLER_82_377 ();
 decap_12 FILLER_82_389 ();
 decap_12 FILLER_82_401 ();
 fill_4 FILLER_82_413 ();
 fill_2 FILLER_82_417 ();
 fill_1 FILLER_82_419 ();
 decap_12 FILLER_82_421 ();
 decap_12 FILLER_82_433 ();
 decap_12 FILLER_82_445 ();
 decap_12 FILLER_82_457 ();
 fill_4 FILLER_82_469 ();
 fill_2 FILLER_82_473 ();
 fill_1 FILLER_82_475 ();
 decap_12 FILLER_82_477 ();
 decap_12 FILLER_82_489 ();
 decap_12 FILLER_82_501 ();
 decap_12 FILLER_82_513 ();
 fill_4 FILLER_82_525 ();
 fill_2 FILLER_82_529 ();
 fill_1 FILLER_82_531 ();
 decap_12 FILLER_82_533 ();
 decap_12 FILLER_82_545 ();
 decap_12 FILLER_82_557 ();
 decap_12 FILLER_82_569 ();
 fill_4 FILLER_82_581 ();
 fill_2 FILLER_82_585 ();
 fill_1 FILLER_82_587 ();
 decap_12 FILLER_82_589 ();
 decap_12 FILLER_82_601 ();
 decap_12 FILLER_82_613 ();
 decap_12 FILLER_83_3 ();
 decap_12 FILLER_83_15 ();
 decap_12 FILLER_83_27 ();
 decap_12 FILLER_83_39 ();
 fill_4 FILLER_83_51 ();
 fill_1 FILLER_83_55 ();
 decap_12 FILLER_83_57 ();
 decap_12 FILLER_83_69 ();
 decap_12 FILLER_83_81 ();
 decap_12 FILLER_83_93 ();
 fill_4 FILLER_83_105 ();
 fill_2 FILLER_83_109 ();
 fill_1 FILLER_83_111 ();
 decap_12 FILLER_83_113 ();
 decap_12 FILLER_83_125 ();
 decap_12 FILLER_83_137 ();
 decap_12 FILLER_83_149 ();
 fill_4 FILLER_83_161 ();
 fill_2 FILLER_83_165 ();
 fill_1 FILLER_83_167 ();
 decap_12 FILLER_83_169 ();
 decap_12 FILLER_83_181 ();
 decap_12 FILLER_83_193 ();
 decap_12 FILLER_83_205 ();
 fill_4 FILLER_83_217 ();
 fill_2 FILLER_83_221 ();
 fill_1 FILLER_83_223 ();
 decap_12 FILLER_83_225 ();
 decap_12 FILLER_83_237 ();
 decap_12 FILLER_83_249 ();
 decap_12 FILLER_83_261 ();
 fill_4 FILLER_83_273 ();
 fill_2 FILLER_83_277 ();
 fill_1 FILLER_83_279 ();
 decap_12 FILLER_83_281 ();
 decap_12 FILLER_83_293 ();
 decap_12 FILLER_83_305 ();
 decap_12 FILLER_83_317 ();
 fill_4 FILLER_83_329 ();
 fill_2 FILLER_83_333 ();
 fill_1 FILLER_83_335 ();
 decap_12 FILLER_83_337 ();
 decap_12 FILLER_83_349 ();
 decap_12 FILLER_83_361 ();
 decap_12 FILLER_83_373 ();
 fill_4 FILLER_83_385 ();
 fill_2 FILLER_83_389 ();
 fill_1 FILLER_83_391 ();
 decap_12 FILLER_83_393 ();
 decap_12 FILLER_83_405 ();
 decap_12 FILLER_83_417 ();
 decap_12 FILLER_83_429 ();
 fill_4 FILLER_83_441 ();
 fill_2 FILLER_83_445 ();
 fill_1 FILLER_83_447 ();
 decap_12 FILLER_83_449 ();
 decap_12 FILLER_83_461 ();
 decap_12 FILLER_83_473 ();
 decap_12 FILLER_83_485 ();
 fill_4 FILLER_83_497 ();
 fill_2 FILLER_83_501 ();
 fill_1 FILLER_83_503 ();
 decap_12 FILLER_83_505 ();
 decap_12 FILLER_83_517 ();
 decap_12 FILLER_83_529 ();
 decap_12 FILLER_83_541 ();
 fill_4 FILLER_83_553 ();
 fill_2 FILLER_83_557 ();
 fill_1 FILLER_83_559 ();
 decap_12 FILLER_83_561 ();
 decap_12 FILLER_83_573 ();
 decap_12 FILLER_83_585 ();
 decap_12 FILLER_83_597 ();
 fill_4 FILLER_83_609 ();
 fill_2 FILLER_83_613 ();
 fill_1 FILLER_83_615 ();
 fill_8 FILLER_83_617 ();
 decap_12 FILLER_84_3 ();
 decap_12 FILLER_84_15 ();
 fill_1 FILLER_84_27 ();
 decap_12 FILLER_84_29 ();
 decap_12 FILLER_84_41 ();
 decap_12 FILLER_84_53 ();
 decap_12 FILLER_84_65 ();
 fill_4 FILLER_84_77 ();
 fill_2 FILLER_84_81 ();
 fill_1 FILLER_84_83 ();
 decap_12 FILLER_84_85 ();
 decap_12 FILLER_84_97 ();
 decap_12 FILLER_84_109 ();
 decap_12 FILLER_84_121 ();
 fill_4 FILLER_84_133 ();
 fill_2 FILLER_84_137 ();
 fill_1 FILLER_84_139 ();
 decap_12 FILLER_84_141 ();
 decap_12 FILLER_84_153 ();
 decap_12 FILLER_84_165 ();
 decap_12 FILLER_84_177 ();
 fill_4 FILLER_84_189 ();
 fill_2 FILLER_84_193 ();
 fill_1 FILLER_84_195 ();
 decap_12 FILLER_84_197 ();
 decap_12 FILLER_84_209 ();
 decap_12 FILLER_84_221 ();
 decap_12 FILLER_84_233 ();
 fill_4 FILLER_84_245 ();
 fill_2 FILLER_84_249 ();
 fill_1 FILLER_84_251 ();
 decap_12 FILLER_84_253 ();
 decap_12 FILLER_84_265 ();
 decap_12 FILLER_84_277 ();
 decap_12 FILLER_84_289 ();
 fill_4 FILLER_84_301 ();
 fill_2 FILLER_84_305 ();
 fill_1 FILLER_84_307 ();
 decap_12 FILLER_84_309 ();
 decap_12 FILLER_84_321 ();
 decap_12 FILLER_84_333 ();
 decap_12 FILLER_84_345 ();
 fill_4 FILLER_84_357 ();
 fill_2 FILLER_84_361 ();
 fill_1 FILLER_84_363 ();
 decap_12 FILLER_84_365 ();
 decap_12 FILLER_84_377 ();
 decap_12 FILLER_84_389 ();
 decap_12 FILLER_84_401 ();
 fill_4 FILLER_84_413 ();
 fill_2 FILLER_84_417 ();
 fill_1 FILLER_84_419 ();
 decap_12 FILLER_84_421 ();
 decap_12 FILLER_84_433 ();
 decap_12 FILLER_84_445 ();
 decap_12 FILLER_84_457 ();
 fill_4 FILLER_84_469 ();
 fill_2 FILLER_84_473 ();
 fill_1 FILLER_84_475 ();
 decap_12 FILLER_84_477 ();
 decap_12 FILLER_84_489 ();
 decap_12 FILLER_84_501 ();
 decap_12 FILLER_84_513 ();
 fill_4 FILLER_84_525 ();
 fill_2 FILLER_84_529 ();
 fill_1 FILLER_84_531 ();
 decap_12 FILLER_84_533 ();
 decap_12 FILLER_84_545 ();
 decap_12 FILLER_84_557 ();
 decap_12 FILLER_84_569 ();
 fill_4 FILLER_84_581 ();
 fill_2 FILLER_84_585 ();
 fill_1 FILLER_84_587 ();
 decap_12 FILLER_84_589 ();
 decap_12 FILLER_84_601 ();
 decap_12 FILLER_84_613 ();
 decap_12 FILLER_85_3 ();
 decap_12 FILLER_85_15 ();
 decap_12 FILLER_85_27 ();
 decap_12 FILLER_85_39 ();
 fill_4 FILLER_85_51 ();
 fill_1 FILLER_85_55 ();
 decap_12 FILLER_85_57 ();
 decap_12 FILLER_85_69 ();
 decap_12 FILLER_85_81 ();
 decap_12 FILLER_85_93 ();
 fill_4 FILLER_85_105 ();
 fill_2 FILLER_85_109 ();
 fill_1 FILLER_85_111 ();
 decap_12 FILLER_85_113 ();
 decap_12 FILLER_85_125 ();
 decap_12 FILLER_85_137 ();
 decap_12 FILLER_85_149 ();
 fill_4 FILLER_85_161 ();
 fill_2 FILLER_85_165 ();
 fill_1 FILLER_85_167 ();
 decap_12 FILLER_85_169 ();
 decap_12 FILLER_85_181 ();
 decap_12 FILLER_85_193 ();
 decap_12 FILLER_85_205 ();
 fill_4 FILLER_85_217 ();
 fill_2 FILLER_85_221 ();
 fill_1 FILLER_85_223 ();
 decap_12 FILLER_85_225 ();
 decap_12 FILLER_85_237 ();
 decap_12 FILLER_85_249 ();
 decap_12 FILLER_85_261 ();
 fill_4 FILLER_85_273 ();
 fill_2 FILLER_85_277 ();
 fill_1 FILLER_85_279 ();
 decap_12 FILLER_85_281 ();
 decap_12 FILLER_85_293 ();
 decap_12 FILLER_85_305 ();
 decap_12 FILLER_85_317 ();
 fill_4 FILLER_85_329 ();
 fill_2 FILLER_85_333 ();
 fill_1 FILLER_85_335 ();
 decap_12 FILLER_85_337 ();
 decap_12 FILLER_85_349 ();
 decap_12 FILLER_85_361 ();
 decap_12 FILLER_85_373 ();
 fill_4 FILLER_85_385 ();
 fill_2 FILLER_85_389 ();
 fill_1 FILLER_85_391 ();
 decap_12 FILLER_85_393 ();
 decap_12 FILLER_85_405 ();
 decap_12 FILLER_85_417 ();
 decap_12 FILLER_85_429 ();
 fill_4 FILLER_85_441 ();
 fill_2 FILLER_85_445 ();
 fill_1 FILLER_85_447 ();
 decap_12 FILLER_85_449 ();
 decap_12 FILLER_85_461 ();
 decap_12 FILLER_85_473 ();
 decap_12 FILLER_85_485 ();
 fill_4 FILLER_85_497 ();
 fill_2 FILLER_85_501 ();
 fill_1 FILLER_85_503 ();
 decap_12 FILLER_85_505 ();
 decap_12 FILLER_85_517 ();
 decap_12 FILLER_85_529 ();
 decap_12 FILLER_85_541 ();
 fill_4 FILLER_85_553 ();
 fill_2 FILLER_85_557 ();
 fill_1 FILLER_85_559 ();
 decap_12 FILLER_85_561 ();
 decap_12 FILLER_85_573 ();
 decap_12 FILLER_85_585 ();
 decap_12 FILLER_85_597 ();
 fill_4 FILLER_85_609 ();
 fill_2 FILLER_85_613 ();
 fill_1 FILLER_85_615 ();
 fill_8 FILLER_85_617 ();
 decap_12 FILLER_86_3 ();
 decap_12 FILLER_86_15 ();
 fill_1 FILLER_86_27 ();
 decap_12 FILLER_86_29 ();
 decap_12 FILLER_86_41 ();
 decap_12 FILLER_86_53 ();
 decap_12 FILLER_86_65 ();
 fill_4 FILLER_86_77 ();
 fill_2 FILLER_86_81 ();
 fill_1 FILLER_86_83 ();
 decap_12 FILLER_86_85 ();
 decap_12 FILLER_86_97 ();
 decap_12 FILLER_86_109 ();
 decap_12 FILLER_86_121 ();
 fill_4 FILLER_86_133 ();
 fill_2 FILLER_86_137 ();
 fill_1 FILLER_86_139 ();
 decap_12 FILLER_86_141 ();
 decap_12 FILLER_86_153 ();
 decap_12 FILLER_86_165 ();
 decap_12 FILLER_86_177 ();
 fill_4 FILLER_86_189 ();
 fill_2 FILLER_86_193 ();
 fill_1 FILLER_86_195 ();
 decap_12 FILLER_86_197 ();
 decap_12 FILLER_86_209 ();
 decap_12 FILLER_86_221 ();
 decap_12 FILLER_86_233 ();
 fill_4 FILLER_86_245 ();
 fill_2 FILLER_86_249 ();
 fill_1 FILLER_86_251 ();
 decap_12 FILLER_86_253 ();
 decap_12 FILLER_86_265 ();
 decap_12 FILLER_86_277 ();
 decap_12 FILLER_86_289 ();
 fill_4 FILLER_86_301 ();
 fill_2 FILLER_86_305 ();
 fill_1 FILLER_86_307 ();
 decap_12 FILLER_86_309 ();
 decap_12 FILLER_86_321 ();
 decap_12 FILLER_86_333 ();
 decap_12 FILLER_86_345 ();
 fill_4 FILLER_86_357 ();
 fill_2 FILLER_86_361 ();
 fill_1 FILLER_86_363 ();
 decap_12 FILLER_86_365 ();
 decap_12 FILLER_86_377 ();
 decap_12 FILLER_86_389 ();
 decap_12 FILLER_86_401 ();
 fill_4 FILLER_86_413 ();
 fill_2 FILLER_86_417 ();
 fill_1 FILLER_86_419 ();
 decap_12 FILLER_86_421 ();
 decap_12 FILLER_86_433 ();
 decap_12 FILLER_86_445 ();
 decap_12 FILLER_86_457 ();
 fill_4 FILLER_86_469 ();
 fill_2 FILLER_86_473 ();
 fill_1 FILLER_86_475 ();
 decap_12 FILLER_86_477 ();
 decap_12 FILLER_86_489 ();
 decap_12 FILLER_86_501 ();
 decap_12 FILLER_86_513 ();
 fill_4 FILLER_86_525 ();
 fill_2 FILLER_86_529 ();
 fill_1 FILLER_86_531 ();
 decap_12 FILLER_86_533 ();
 decap_12 FILLER_86_545 ();
 decap_12 FILLER_86_557 ();
 decap_12 FILLER_86_569 ();
 fill_4 FILLER_86_581 ();
 fill_2 FILLER_86_585 ();
 fill_1 FILLER_86_587 ();
 decap_12 FILLER_86_589 ();
 decap_12 FILLER_86_601 ();
 decap_12 FILLER_86_613 ();
 decap_12 FILLER_87_3 ();
 decap_12 FILLER_87_15 ();
 decap_12 FILLER_87_27 ();
 decap_12 FILLER_87_39 ();
 fill_4 FILLER_87_51 ();
 fill_1 FILLER_87_55 ();
 decap_12 FILLER_87_57 ();
 decap_12 FILLER_87_69 ();
 decap_12 FILLER_87_81 ();
 decap_12 FILLER_87_93 ();
 fill_4 FILLER_87_105 ();
 fill_2 FILLER_87_109 ();
 fill_1 FILLER_87_111 ();
 decap_12 FILLER_87_113 ();
 decap_12 FILLER_87_125 ();
 decap_12 FILLER_87_137 ();
 decap_12 FILLER_87_149 ();
 fill_4 FILLER_87_161 ();
 fill_2 FILLER_87_165 ();
 fill_1 FILLER_87_167 ();
 decap_12 FILLER_87_169 ();
 decap_12 FILLER_87_181 ();
 decap_12 FILLER_87_193 ();
 decap_12 FILLER_87_205 ();
 fill_4 FILLER_87_217 ();
 fill_2 FILLER_87_221 ();
 fill_1 FILLER_87_223 ();
 decap_12 FILLER_87_225 ();
 decap_12 FILLER_87_237 ();
 decap_12 FILLER_87_249 ();
 decap_12 FILLER_87_261 ();
 fill_4 FILLER_87_273 ();
 fill_2 FILLER_87_277 ();
 fill_1 FILLER_87_279 ();
 decap_12 FILLER_87_281 ();
 decap_12 FILLER_87_293 ();
 decap_12 FILLER_87_305 ();
 decap_12 FILLER_87_317 ();
 fill_4 FILLER_87_329 ();
 fill_2 FILLER_87_333 ();
 fill_1 FILLER_87_335 ();
 decap_12 FILLER_87_337 ();
 decap_12 FILLER_87_349 ();
 decap_12 FILLER_87_361 ();
 decap_12 FILLER_87_373 ();
 fill_4 FILLER_87_385 ();
 fill_2 FILLER_87_389 ();
 fill_1 FILLER_87_391 ();
 decap_12 FILLER_87_393 ();
 decap_12 FILLER_87_405 ();
 decap_12 FILLER_87_417 ();
 decap_12 FILLER_87_429 ();
 fill_4 FILLER_87_441 ();
 fill_2 FILLER_87_445 ();
 fill_1 FILLER_87_447 ();
 decap_12 FILLER_87_449 ();
 decap_12 FILLER_87_461 ();
 decap_12 FILLER_87_473 ();
 decap_12 FILLER_87_485 ();
 fill_4 FILLER_87_497 ();
 fill_2 FILLER_87_501 ();
 fill_1 FILLER_87_503 ();
 decap_12 FILLER_87_505 ();
 decap_12 FILLER_87_517 ();
 decap_12 FILLER_87_529 ();
 decap_12 FILLER_87_541 ();
 fill_4 FILLER_87_553 ();
 fill_2 FILLER_87_557 ();
 fill_1 FILLER_87_559 ();
 decap_12 FILLER_87_561 ();
 decap_12 FILLER_87_573 ();
 decap_12 FILLER_87_585 ();
 decap_12 FILLER_87_597 ();
 fill_4 FILLER_87_609 ();
 fill_2 FILLER_87_613 ();
 fill_1 FILLER_87_615 ();
 fill_8 FILLER_87_617 ();
 decap_12 FILLER_88_3 ();
 decap_12 FILLER_88_15 ();
 fill_1 FILLER_88_27 ();
 decap_12 FILLER_88_29 ();
 decap_12 FILLER_88_41 ();
 decap_12 FILLER_88_53 ();
 decap_12 FILLER_88_65 ();
 fill_4 FILLER_88_77 ();
 fill_2 FILLER_88_81 ();
 fill_1 FILLER_88_83 ();
 decap_12 FILLER_88_85 ();
 decap_12 FILLER_88_97 ();
 decap_12 FILLER_88_109 ();
 decap_12 FILLER_88_121 ();
 fill_4 FILLER_88_133 ();
 fill_2 FILLER_88_137 ();
 fill_1 FILLER_88_139 ();
 decap_12 FILLER_88_141 ();
 decap_12 FILLER_88_153 ();
 decap_12 FILLER_88_165 ();
 decap_12 FILLER_88_177 ();
 fill_4 FILLER_88_189 ();
 fill_2 FILLER_88_193 ();
 fill_1 FILLER_88_195 ();
 decap_12 FILLER_88_197 ();
 decap_12 FILLER_88_209 ();
 decap_12 FILLER_88_221 ();
 decap_12 FILLER_88_233 ();
 fill_4 FILLER_88_245 ();
 fill_2 FILLER_88_249 ();
 fill_1 FILLER_88_251 ();
 decap_12 FILLER_88_253 ();
 decap_12 FILLER_88_265 ();
 decap_12 FILLER_88_277 ();
 decap_12 FILLER_88_289 ();
 fill_4 FILLER_88_301 ();
 fill_2 FILLER_88_305 ();
 fill_1 FILLER_88_307 ();
 decap_12 FILLER_88_309 ();
 decap_12 FILLER_88_321 ();
 decap_12 FILLER_88_333 ();
 decap_12 FILLER_88_345 ();
 fill_4 FILLER_88_357 ();
 fill_2 FILLER_88_361 ();
 fill_1 FILLER_88_363 ();
 decap_12 FILLER_88_365 ();
 decap_12 FILLER_88_377 ();
 decap_12 FILLER_88_389 ();
 decap_12 FILLER_88_401 ();
 fill_4 FILLER_88_413 ();
 fill_2 FILLER_88_417 ();
 fill_1 FILLER_88_419 ();
 decap_12 FILLER_88_421 ();
 decap_12 FILLER_88_433 ();
 decap_12 FILLER_88_445 ();
 decap_12 FILLER_88_457 ();
 fill_4 FILLER_88_469 ();
 fill_2 FILLER_88_473 ();
 fill_1 FILLER_88_475 ();
 decap_12 FILLER_88_477 ();
 decap_12 FILLER_88_489 ();
 decap_12 FILLER_88_501 ();
 decap_12 FILLER_88_513 ();
 fill_4 FILLER_88_525 ();
 fill_2 FILLER_88_529 ();
 fill_1 FILLER_88_531 ();
 decap_12 FILLER_88_533 ();
 decap_12 FILLER_88_545 ();
 decap_12 FILLER_88_557 ();
 decap_12 FILLER_88_569 ();
 fill_4 FILLER_88_581 ();
 fill_2 FILLER_88_585 ();
 fill_1 FILLER_88_587 ();
 decap_12 FILLER_88_589 ();
 decap_12 FILLER_88_601 ();
 decap_12 FILLER_88_613 ();
 decap_12 FILLER_89_3 ();
 decap_12 FILLER_89_15 ();
 decap_12 FILLER_89_27 ();
 decap_12 FILLER_89_39 ();
 fill_4 FILLER_89_51 ();
 fill_1 FILLER_89_55 ();
 decap_12 FILLER_89_57 ();
 decap_12 FILLER_89_69 ();
 decap_12 FILLER_89_81 ();
 decap_12 FILLER_89_93 ();
 fill_4 FILLER_89_105 ();
 fill_2 FILLER_89_109 ();
 fill_1 FILLER_89_111 ();
 decap_12 FILLER_89_113 ();
 decap_12 FILLER_89_125 ();
 decap_12 FILLER_89_137 ();
 decap_12 FILLER_89_149 ();
 fill_4 FILLER_89_161 ();
 fill_2 FILLER_89_165 ();
 fill_1 FILLER_89_167 ();
 decap_12 FILLER_89_169 ();
 decap_12 FILLER_89_181 ();
 decap_12 FILLER_89_193 ();
 decap_12 FILLER_89_205 ();
 fill_4 FILLER_89_217 ();
 fill_2 FILLER_89_221 ();
 fill_1 FILLER_89_223 ();
 decap_12 FILLER_89_225 ();
 decap_12 FILLER_89_237 ();
 decap_12 FILLER_89_249 ();
 decap_12 FILLER_89_261 ();
 fill_4 FILLER_89_273 ();
 fill_2 FILLER_89_277 ();
 fill_1 FILLER_89_279 ();
 decap_12 FILLER_89_281 ();
 decap_12 FILLER_89_293 ();
 decap_12 FILLER_89_305 ();
 decap_12 FILLER_89_317 ();
 fill_4 FILLER_89_329 ();
 fill_2 FILLER_89_333 ();
 fill_1 FILLER_89_335 ();
 decap_12 FILLER_89_337 ();
 decap_12 FILLER_89_349 ();
 decap_12 FILLER_89_361 ();
 decap_12 FILLER_89_373 ();
 fill_4 FILLER_89_385 ();
 fill_2 FILLER_89_389 ();
 fill_1 FILLER_89_391 ();
 decap_12 FILLER_89_393 ();
 decap_12 FILLER_89_405 ();
 decap_12 FILLER_89_417 ();
 decap_12 FILLER_89_429 ();
 fill_4 FILLER_89_441 ();
 fill_2 FILLER_89_445 ();
 fill_1 FILLER_89_447 ();
 decap_12 FILLER_89_449 ();
 decap_12 FILLER_89_461 ();
 decap_12 FILLER_89_473 ();
 decap_12 FILLER_89_485 ();
 fill_4 FILLER_89_497 ();
 fill_2 FILLER_89_501 ();
 fill_1 FILLER_89_503 ();
 decap_12 FILLER_89_505 ();
 decap_12 FILLER_89_517 ();
 decap_12 FILLER_89_529 ();
 decap_12 FILLER_89_541 ();
 fill_4 FILLER_89_553 ();
 fill_2 FILLER_89_557 ();
 fill_1 FILLER_89_559 ();
 decap_12 FILLER_89_561 ();
 decap_12 FILLER_89_573 ();
 decap_12 FILLER_89_585 ();
 decap_12 FILLER_89_597 ();
 fill_4 FILLER_89_609 ();
 fill_2 FILLER_89_613 ();
 fill_1 FILLER_89_615 ();
 fill_8 FILLER_89_617 ();
 decap_12 FILLER_90_3 ();
 decap_12 FILLER_90_15 ();
 fill_1 FILLER_90_27 ();
 decap_12 FILLER_90_29 ();
 decap_12 FILLER_90_41 ();
 decap_12 FILLER_90_53 ();
 decap_12 FILLER_90_65 ();
 fill_4 FILLER_90_77 ();
 fill_2 FILLER_90_81 ();
 fill_1 FILLER_90_83 ();
 decap_12 FILLER_90_85 ();
 decap_12 FILLER_90_97 ();
 decap_12 FILLER_90_109 ();
 decap_12 FILLER_90_121 ();
 fill_4 FILLER_90_133 ();
 fill_2 FILLER_90_137 ();
 fill_1 FILLER_90_139 ();
 decap_12 FILLER_90_141 ();
 decap_12 FILLER_90_153 ();
 decap_12 FILLER_90_165 ();
 decap_12 FILLER_90_177 ();
 fill_4 FILLER_90_189 ();
 fill_2 FILLER_90_193 ();
 fill_1 FILLER_90_195 ();
 decap_12 FILLER_90_197 ();
 decap_12 FILLER_90_209 ();
 decap_12 FILLER_90_221 ();
 decap_12 FILLER_90_233 ();
 fill_4 FILLER_90_245 ();
 fill_2 FILLER_90_249 ();
 fill_1 FILLER_90_251 ();
 decap_12 FILLER_90_253 ();
 decap_12 FILLER_90_265 ();
 decap_12 FILLER_90_277 ();
 decap_12 FILLER_90_289 ();
 fill_4 FILLER_90_301 ();
 fill_2 FILLER_90_305 ();
 fill_1 FILLER_90_307 ();
 decap_12 FILLER_90_309 ();
 decap_12 FILLER_90_321 ();
 decap_12 FILLER_90_333 ();
 decap_12 FILLER_90_345 ();
 fill_4 FILLER_90_357 ();
 fill_2 FILLER_90_361 ();
 fill_1 FILLER_90_363 ();
 decap_12 FILLER_90_365 ();
 decap_12 FILLER_90_377 ();
 decap_12 FILLER_90_389 ();
 decap_12 FILLER_90_401 ();
 fill_4 FILLER_90_413 ();
 fill_2 FILLER_90_417 ();
 fill_1 FILLER_90_419 ();
 decap_12 FILLER_90_421 ();
 decap_12 FILLER_90_433 ();
 decap_12 FILLER_90_445 ();
 decap_12 FILLER_90_457 ();
 fill_4 FILLER_90_469 ();
 fill_2 FILLER_90_473 ();
 fill_1 FILLER_90_475 ();
 decap_12 FILLER_90_477 ();
 decap_12 FILLER_90_489 ();
 decap_12 FILLER_90_501 ();
 decap_12 FILLER_90_513 ();
 fill_4 FILLER_90_525 ();
 fill_2 FILLER_90_529 ();
 fill_1 FILLER_90_531 ();
 decap_12 FILLER_90_533 ();
 decap_12 FILLER_90_545 ();
 decap_12 FILLER_90_557 ();
 decap_12 FILLER_90_569 ();
 fill_4 FILLER_90_581 ();
 fill_2 FILLER_90_585 ();
 fill_1 FILLER_90_587 ();
 decap_12 FILLER_90_589 ();
 decap_12 FILLER_90_601 ();
 decap_12 FILLER_90_613 ();
 decap_12 FILLER_91_3 ();
 decap_12 FILLER_91_15 ();
 decap_12 FILLER_91_27 ();
 decap_12 FILLER_91_39 ();
 fill_4 FILLER_91_51 ();
 fill_1 FILLER_91_55 ();
 decap_12 FILLER_91_57 ();
 decap_12 FILLER_91_69 ();
 decap_12 FILLER_91_81 ();
 decap_12 FILLER_91_93 ();
 fill_4 FILLER_91_105 ();
 fill_2 FILLER_91_109 ();
 fill_1 FILLER_91_111 ();
 decap_12 FILLER_91_113 ();
 decap_12 FILLER_91_125 ();
 decap_12 FILLER_91_137 ();
 decap_12 FILLER_91_149 ();
 fill_4 FILLER_91_161 ();
 fill_2 FILLER_91_165 ();
 fill_1 FILLER_91_167 ();
 decap_12 FILLER_91_169 ();
 decap_12 FILLER_91_181 ();
 decap_12 FILLER_91_193 ();
 decap_12 FILLER_91_205 ();
 fill_4 FILLER_91_217 ();
 fill_2 FILLER_91_221 ();
 fill_1 FILLER_91_223 ();
 decap_12 FILLER_91_225 ();
 decap_12 FILLER_91_237 ();
 decap_12 FILLER_91_249 ();
 decap_12 FILLER_91_261 ();
 fill_4 FILLER_91_273 ();
 fill_2 FILLER_91_277 ();
 fill_1 FILLER_91_279 ();
 decap_12 FILLER_91_281 ();
 decap_12 FILLER_91_293 ();
 decap_12 FILLER_91_305 ();
 decap_12 FILLER_91_317 ();
 fill_4 FILLER_91_329 ();
 fill_2 FILLER_91_333 ();
 fill_1 FILLER_91_335 ();
 decap_12 FILLER_91_337 ();
 decap_12 FILLER_91_349 ();
 decap_12 FILLER_91_361 ();
 decap_12 FILLER_91_373 ();
 fill_4 FILLER_91_385 ();
 fill_2 FILLER_91_389 ();
 fill_1 FILLER_91_391 ();
 decap_12 FILLER_91_393 ();
 decap_12 FILLER_91_405 ();
 decap_12 FILLER_91_417 ();
 decap_12 FILLER_91_429 ();
 fill_4 FILLER_91_441 ();
 fill_2 FILLER_91_445 ();
 fill_1 FILLER_91_447 ();
 decap_12 FILLER_91_449 ();
 decap_12 FILLER_91_461 ();
 decap_12 FILLER_91_473 ();
 decap_12 FILLER_91_485 ();
 fill_4 FILLER_91_497 ();
 fill_2 FILLER_91_501 ();
 fill_1 FILLER_91_503 ();
 decap_12 FILLER_91_505 ();
 decap_12 FILLER_91_517 ();
 decap_12 FILLER_91_529 ();
 decap_12 FILLER_91_541 ();
 fill_4 FILLER_91_553 ();
 fill_2 FILLER_91_557 ();
 fill_1 FILLER_91_559 ();
 decap_12 FILLER_91_561 ();
 decap_12 FILLER_91_573 ();
 decap_12 FILLER_91_585 ();
 decap_12 FILLER_91_597 ();
 fill_4 FILLER_91_609 ();
 fill_2 FILLER_91_613 ();
 fill_1 FILLER_91_615 ();
 fill_8 FILLER_91_617 ();
 decap_12 FILLER_92_3 ();
 decap_12 FILLER_92_15 ();
 fill_1 FILLER_92_27 ();
 decap_12 FILLER_92_29 ();
 decap_12 FILLER_92_41 ();
 decap_12 FILLER_92_53 ();
 decap_12 FILLER_92_65 ();
 fill_4 FILLER_92_77 ();
 fill_2 FILLER_92_81 ();
 fill_1 FILLER_92_83 ();
 decap_12 FILLER_92_85 ();
 decap_12 FILLER_92_97 ();
 decap_12 FILLER_92_109 ();
 decap_12 FILLER_92_121 ();
 fill_4 FILLER_92_133 ();
 fill_2 FILLER_92_137 ();
 fill_1 FILLER_92_139 ();
 decap_12 FILLER_92_141 ();
 decap_12 FILLER_92_153 ();
 decap_12 FILLER_92_165 ();
 decap_12 FILLER_92_177 ();
 fill_4 FILLER_92_189 ();
 fill_2 FILLER_92_193 ();
 fill_1 FILLER_92_195 ();
 decap_12 FILLER_92_197 ();
 decap_12 FILLER_92_209 ();
 decap_12 FILLER_92_221 ();
 decap_12 FILLER_92_233 ();
 fill_4 FILLER_92_245 ();
 fill_2 FILLER_92_249 ();
 fill_1 FILLER_92_251 ();
 decap_12 FILLER_92_253 ();
 decap_12 FILLER_92_265 ();
 decap_12 FILLER_92_277 ();
 decap_12 FILLER_92_289 ();
 fill_4 FILLER_92_301 ();
 fill_2 FILLER_92_305 ();
 fill_1 FILLER_92_307 ();
 decap_12 FILLER_92_309 ();
 decap_12 FILLER_92_321 ();
 decap_12 FILLER_92_333 ();
 decap_12 FILLER_92_345 ();
 fill_4 FILLER_92_357 ();
 fill_2 FILLER_92_361 ();
 fill_1 FILLER_92_363 ();
 decap_12 FILLER_92_365 ();
 decap_12 FILLER_92_377 ();
 decap_12 FILLER_92_389 ();
 decap_12 FILLER_92_401 ();
 fill_4 FILLER_92_413 ();
 fill_2 FILLER_92_417 ();
 fill_1 FILLER_92_419 ();
 decap_12 FILLER_92_421 ();
 decap_12 FILLER_92_433 ();
 decap_12 FILLER_92_445 ();
 decap_12 FILLER_92_457 ();
 fill_4 FILLER_92_469 ();
 fill_2 FILLER_92_473 ();
 fill_1 FILLER_92_475 ();
 decap_12 FILLER_92_477 ();
 decap_12 FILLER_92_489 ();
 decap_12 FILLER_92_501 ();
 decap_12 FILLER_92_513 ();
 fill_4 FILLER_92_525 ();
 fill_2 FILLER_92_529 ();
 fill_1 FILLER_92_531 ();
 decap_12 FILLER_92_533 ();
 decap_12 FILLER_92_545 ();
 decap_12 FILLER_92_557 ();
 decap_12 FILLER_92_569 ();
 fill_4 FILLER_92_581 ();
 fill_2 FILLER_92_585 ();
 fill_1 FILLER_92_587 ();
 decap_12 FILLER_92_589 ();
 decap_12 FILLER_92_601 ();
 decap_12 FILLER_92_613 ();
 decap_12 FILLER_93_3 ();
 decap_12 FILLER_93_15 ();
 decap_12 FILLER_93_27 ();
 decap_12 FILLER_93_39 ();
 fill_4 FILLER_93_51 ();
 fill_1 FILLER_93_55 ();
 decap_12 FILLER_93_57 ();
 decap_12 FILLER_93_69 ();
 decap_12 FILLER_93_81 ();
 decap_12 FILLER_93_93 ();
 fill_4 FILLER_93_105 ();
 fill_2 FILLER_93_109 ();
 fill_1 FILLER_93_111 ();
 decap_12 FILLER_93_113 ();
 decap_12 FILLER_93_125 ();
 decap_12 FILLER_93_137 ();
 decap_12 FILLER_93_149 ();
 fill_4 FILLER_93_161 ();
 fill_2 FILLER_93_165 ();
 fill_1 FILLER_93_167 ();
 decap_12 FILLER_93_169 ();
 decap_12 FILLER_93_181 ();
 decap_12 FILLER_93_193 ();
 decap_12 FILLER_93_205 ();
 fill_4 FILLER_93_217 ();
 fill_2 FILLER_93_221 ();
 fill_1 FILLER_93_223 ();
 decap_12 FILLER_93_225 ();
 decap_12 FILLER_93_237 ();
 decap_12 FILLER_93_249 ();
 decap_12 FILLER_93_261 ();
 fill_4 FILLER_93_273 ();
 fill_2 FILLER_93_277 ();
 fill_1 FILLER_93_279 ();
 decap_12 FILLER_93_281 ();
 decap_12 FILLER_93_293 ();
 decap_12 FILLER_93_305 ();
 decap_12 FILLER_93_317 ();
 fill_4 FILLER_93_329 ();
 fill_2 FILLER_93_333 ();
 fill_1 FILLER_93_335 ();
 decap_12 FILLER_93_337 ();
 decap_12 FILLER_93_349 ();
 decap_12 FILLER_93_361 ();
 decap_12 FILLER_93_373 ();
 fill_4 FILLER_93_385 ();
 fill_2 FILLER_93_389 ();
 fill_1 FILLER_93_391 ();
 decap_12 FILLER_93_393 ();
 decap_12 FILLER_93_405 ();
 decap_12 FILLER_93_417 ();
 decap_12 FILLER_93_429 ();
 fill_4 FILLER_93_441 ();
 fill_2 FILLER_93_445 ();
 fill_1 FILLER_93_447 ();
 decap_12 FILLER_93_449 ();
 decap_12 FILLER_93_461 ();
 decap_12 FILLER_93_473 ();
 decap_12 FILLER_93_485 ();
 fill_4 FILLER_93_497 ();
 fill_2 FILLER_93_501 ();
 fill_1 FILLER_93_503 ();
 decap_12 FILLER_93_505 ();
 decap_12 FILLER_93_517 ();
 decap_12 FILLER_93_529 ();
 decap_12 FILLER_93_541 ();
 fill_4 FILLER_93_553 ();
 fill_2 FILLER_93_557 ();
 fill_1 FILLER_93_559 ();
 decap_12 FILLER_93_561 ();
 decap_12 FILLER_93_573 ();
 decap_12 FILLER_93_585 ();
 decap_12 FILLER_93_597 ();
 fill_4 FILLER_93_609 ();
 fill_2 FILLER_93_613 ();
 fill_1 FILLER_93_615 ();
 fill_8 FILLER_93_617 ();
 decap_12 FILLER_94_3 ();
 decap_12 FILLER_94_15 ();
 fill_1 FILLER_94_27 ();
 decap_12 FILLER_94_29 ();
 decap_12 FILLER_94_41 ();
 decap_12 FILLER_94_53 ();
 decap_12 FILLER_94_65 ();
 fill_4 FILLER_94_77 ();
 fill_2 FILLER_94_81 ();
 fill_1 FILLER_94_83 ();
 decap_12 FILLER_94_85 ();
 decap_12 FILLER_94_97 ();
 decap_12 FILLER_94_109 ();
 decap_12 FILLER_94_121 ();
 fill_4 FILLER_94_133 ();
 fill_2 FILLER_94_137 ();
 fill_1 FILLER_94_139 ();
 decap_12 FILLER_94_141 ();
 decap_12 FILLER_94_153 ();
 decap_12 FILLER_94_165 ();
 decap_12 FILLER_94_177 ();
 fill_4 FILLER_94_189 ();
 fill_2 FILLER_94_193 ();
 fill_1 FILLER_94_195 ();
 decap_12 FILLER_94_197 ();
 decap_12 FILLER_94_209 ();
 decap_12 FILLER_94_221 ();
 decap_12 FILLER_94_233 ();
 fill_4 FILLER_94_245 ();
 fill_2 FILLER_94_249 ();
 fill_1 FILLER_94_251 ();
 decap_12 FILLER_94_253 ();
 decap_12 FILLER_94_265 ();
 decap_12 FILLER_94_277 ();
 decap_12 FILLER_94_289 ();
 fill_4 FILLER_94_301 ();
 fill_2 FILLER_94_305 ();
 fill_1 FILLER_94_307 ();
 decap_12 FILLER_94_309 ();
 decap_12 FILLER_94_321 ();
 decap_12 FILLER_94_333 ();
 decap_12 FILLER_94_345 ();
 fill_4 FILLER_94_357 ();
 fill_2 FILLER_94_361 ();
 fill_1 FILLER_94_363 ();
 decap_12 FILLER_94_365 ();
 decap_12 FILLER_94_377 ();
 decap_12 FILLER_94_389 ();
 decap_12 FILLER_94_401 ();
 fill_4 FILLER_94_413 ();
 fill_2 FILLER_94_417 ();
 fill_1 FILLER_94_419 ();
 decap_12 FILLER_94_421 ();
 decap_12 FILLER_94_433 ();
 decap_12 FILLER_94_445 ();
 decap_12 FILLER_94_457 ();
 fill_4 FILLER_94_469 ();
 fill_2 FILLER_94_473 ();
 fill_1 FILLER_94_475 ();
 decap_12 FILLER_94_477 ();
 decap_12 FILLER_94_489 ();
 decap_12 FILLER_94_501 ();
 decap_12 FILLER_94_513 ();
 fill_4 FILLER_94_525 ();
 fill_2 FILLER_94_529 ();
 fill_1 FILLER_94_531 ();
 decap_12 FILLER_94_533 ();
 decap_12 FILLER_94_545 ();
 decap_12 FILLER_94_557 ();
 decap_12 FILLER_94_569 ();
 fill_4 FILLER_94_581 ();
 fill_2 FILLER_94_585 ();
 fill_1 FILLER_94_587 ();
 decap_12 FILLER_94_589 ();
 decap_12 FILLER_94_601 ();
 decap_12 FILLER_94_613 ();
 decap_12 FILLER_95_3 ();
 decap_12 FILLER_95_15 ();
 decap_12 FILLER_95_27 ();
 decap_12 FILLER_95_39 ();
 fill_4 FILLER_95_51 ();
 fill_1 FILLER_95_55 ();
 decap_12 FILLER_95_57 ();
 decap_12 FILLER_95_69 ();
 decap_12 FILLER_95_81 ();
 decap_12 FILLER_95_93 ();
 fill_4 FILLER_95_105 ();
 fill_2 FILLER_95_109 ();
 fill_1 FILLER_95_111 ();
 decap_12 FILLER_95_113 ();
 decap_12 FILLER_95_125 ();
 decap_12 FILLER_95_137 ();
 decap_12 FILLER_95_149 ();
 fill_4 FILLER_95_161 ();
 fill_2 FILLER_95_165 ();
 fill_1 FILLER_95_167 ();
 decap_12 FILLER_95_169 ();
 decap_12 FILLER_95_181 ();
 decap_12 FILLER_95_193 ();
 decap_12 FILLER_95_205 ();
 fill_4 FILLER_95_217 ();
 fill_2 FILLER_95_221 ();
 fill_1 FILLER_95_223 ();
 decap_12 FILLER_95_225 ();
 decap_12 FILLER_95_237 ();
 decap_12 FILLER_95_249 ();
 decap_12 FILLER_95_261 ();
 fill_4 FILLER_95_273 ();
 fill_2 FILLER_95_277 ();
 fill_1 FILLER_95_279 ();
 decap_12 FILLER_95_281 ();
 decap_12 FILLER_95_293 ();
 decap_12 FILLER_95_305 ();
 decap_12 FILLER_95_317 ();
 fill_4 FILLER_95_329 ();
 fill_2 FILLER_95_333 ();
 fill_1 FILLER_95_335 ();
 decap_12 FILLER_95_337 ();
 decap_12 FILLER_95_349 ();
 decap_12 FILLER_95_361 ();
 decap_12 FILLER_95_373 ();
 fill_4 FILLER_95_385 ();
 fill_2 FILLER_95_389 ();
 fill_1 FILLER_95_391 ();
 decap_12 FILLER_95_393 ();
 decap_12 FILLER_95_405 ();
 decap_12 FILLER_95_417 ();
 decap_12 FILLER_95_429 ();
 fill_4 FILLER_95_441 ();
 fill_2 FILLER_95_445 ();
 fill_1 FILLER_95_447 ();
 decap_12 FILLER_95_449 ();
 decap_12 FILLER_95_461 ();
 decap_12 FILLER_95_473 ();
 decap_12 FILLER_95_485 ();
 fill_4 FILLER_95_497 ();
 fill_2 FILLER_95_501 ();
 fill_1 FILLER_95_503 ();
 decap_12 FILLER_95_505 ();
 decap_12 FILLER_95_517 ();
 decap_12 FILLER_95_529 ();
 decap_12 FILLER_95_541 ();
 fill_4 FILLER_95_553 ();
 fill_2 FILLER_95_557 ();
 fill_1 FILLER_95_559 ();
 decap_12 FILLER_95_561 ();
 decap_12 FILLER_95_573 ();
 decap_12 FILLER_95_585 ();
 decap_12 FILLER_95_597 ();
 fill_4 FILLER_95_609 ();
 fill_2 FILLER_95_613 ();
 fill_1 FILLER_95_615 ();
 fill_8 FILLER_95_617 ();
 decap_12 FILLER_96_3 ();
 decap_12 FILLER_96_15 ();
 fill_1 FILLER_96_27 ();
 decap_12 FILLER_96_29 ();
 decap_12 FILLER_96_41 ();
 decap_12 FILLER_96_53 ();
 decap_12 FILLER_96_65 ();
 fill_4 FILLER_96_77 ();
 fill_2 FILLER_96_81 ();
 fill_1 FILLER_96_83 ();
 decap_12 FILLER_96_85 ();
 decap_12 FILLER_96_97 ();
 decap_12 FILLER_96_109 ();
 decap_12 FILLER_96_121 ();
 fill_4 FILLER_96_133 ();
 fill_2 FILLER_96_137 ();
 fill_1 FILLER_96_139 ();
 decap_12 FILLER_96_141 ();
 decap_12 FILLER_96_153 ();
 decap_12 FILLER_96_165 ();
 decap_12 FILLER_96_177 ();
 fill_4 FILLER_96_189 ();
 fill_2 FILLER_96_193 ();
 fill_1 FILLER_96_195 ();
 decap_12 FILLER_96_197 ();
 decap_12 FILLER_96_209 ();
 decap_12 FILLER_96_221 ();
 decap_12 FILLER_96_233 ();
 fill_4 FILLER_96_245 ();
 fill_2 FILLER_96_249 ();
 fill_1 FILLER_96_251 ();
 decap_12 FILLER_96_253 ();
 decap_12 FILLER_96_265 ();
 decap_12 FILLER_96_277 ();
 decap_12 FILLER_96_289 ();
 fill_4 FILLER_96_301 ();
 fill_2 FILLER_96_305 ();
 fill_1 FILLER_96_307 ();
 decap_12 FILLER_96_309 ();
 decap_12 FILLER_96_321 ();
 decap_12 FILLER_96_333 ();
 decap_12 FILLER_96_345 ();
 fill_4 FILLER_96_357 ();
 fill_2 FILLER_96_361 ();
 fill_1 FILLER_96_363 ();
 decap_12 FILLER_96_365 ();
 decap_12 FILLER_96_377 ();
 decap_12 FILLER_96_389 ();
 decap_12 FILLER_96_401 ();
 fill_4 FILLER_96_413 ();
 fill_2 FILLER_96_417 ();
 fill_1 FILLER_96_419 ();
 decap_12 FILLER_96_421 ();
 decap_12 FILLER_96_433 ();
 decap_12 FILLER_96_445 ();
 decap_12 FILLER_96_457 ();
 fill_4 FILLER_96_469 ();
 fill_2 FILLER_96_473 ();
 fill_1 FILLER_96_475 ();
 decap_12 FILLER_96_477 ();
 decap_12 FILLER_96_489 ();
 decap_12 FILLER_96_501 ();
 decap_12 FILLER_96_513 ();
 fill_4 FILLER_96_525 ();
 fill_2 FILLER_96_529 ();
 fill_1 FILLER_96_531 ();
 decap_12 FILLER_96_533 ();
 decap_12 FILLER_96_545 ();
 decap_12 FILLER_96_557 ();
 decap_12 FILLER_96_569 ();
 fill_4 FILLER_96_581 ();
 fill_2 FILLER_96_585 ();
 fill_1 FILLER_96_587 ();
 decap_12 FILLER_96_589 ();
 decap_12 FILLER_96_601 ();
 decap_12 FILLER_96_613 ();
 decap_12 FILLER_97_3 ();
 decap_12 FILLER_97_15 ();
 decap_12 FILLER_97_27 ();
 decap_12 FILLER_97_39 ();
 fill_4 FILLER_97_51 ();
 fill_1 FILLER_97_55 ();
 decap_12 FILLER_97_57 ();
 decap_12 FILLER_97_69 ();
 decap_12 FILLER_97_81 ();
 decap_12 FILLER_97_93 ();
 fill_4 FILLER_97_105 ();
 fill_2 FILLER_97_109 ();
 fill_1 FILLER_97_111 ();
 decap_12 FILLER_97_113 ();
 decap_12 FILLER_97_125 ();
 decap_12 FILLER_97_137 ();
 decap_12 FILLER_97_149 ();
 fill_4 FILLER_97_161 ();
 fill_2 FILLER_97_165 ();
 fill_1 FILLER_97_167 ();
 decap_12 FILLER_97_169 ();
 decap_12 FILLER_97_181 ();
 decap_12 FILLER_97_193 ();
 decap_12 FILLER_97_205 ();
 fill_4 FILLER_97_217 ();
 fill_2 FILLER_97_221 ();
 fill_1 FILLER_97_223 ();
 decap_12 FILLER_97_225 ();
 decap_12 FILLER_97_237 ();
 decap_12 FILLER_97_249 ();
 decap_12 FILLER_97_261 ();
 fill_4 FILLER_97_273 ();
 fill_2 FILLER_97_277 ();
 fill_1 FILLER_97_279 ();
 decap_12 FILLER_97_281 ();
 decap_12 FILLER_97_293 ();
 decap_12 FILLER_97_305 ();
 decap_12 FILLER_97_317 ();
 fill_4 FILLER_97_329 ();
 fill_2 FILLER_97_333 ();
 fill_1 FILLER_97_335 ();
 decap_12 FILLER_97_337 ();
 decap_12 FILLER_97_349 ();
 decap_12 FILLER_97_361 ();
 decap_12 FILLER_97_373 ();
 fill_4 FILLER_97_385 ();
 fill_2 FILLER_97_389 ();
 fill_1 FILLER_97_391 ();
 decap_12 FILLER_97_393 ();
 decap_12 FILLER_97_405 ();
 decap_12 FILLER_97_417 ();
 decap_12 FILLER_97_429 ();
 fill_4 FILLER_97_441 ();
 fill_2 FILLER_97_445 ();
 fill_1 FILLER_97_447 ();
 decap_12 FILLER_97_449 ();
 decap_12 FILLER_97_461 ();
 decap_12 FILLER_97_473 ();
 decap_12 FILLER_97_485 ();
 fill_4 FILLER_97_497 ();
 fill_2 FILLER_97_501 ();
 fill_1 FILLER_97_503 ();
 decap_12 FILLER_97_505 ();
 decap_12 FILLER_97_517 ();
 decap_12 FILLER_97_529 ();
 decap_12 FILLER_97_541 ();
 fill_4 FILLER_97_553 ();
 fill_2 FILLER_97_557 ();
 fill_1 FILLER_97_559 ();
 decap_12 FILLER_97_561 ();
 decap_12 FILLER_97_573 ();
 decap_12 FILLER_97_585 ();
 decap_12 FILLER_97_597 ();
 fill_4 FILLER_97_609 ();
 fill_2 FILLER_97_613 ();
 fill_1 FILLER_97_615 ();
 fill_8 FILLER_97_617 ();
 decap_12 FILLER_98_3 ();
 decap_12 FILLER_98_15 ();
 fill_1 FILLER_98_27 ();
 decap_12 FILLER_98_29 ();
 decap_12 FILLER_98_41 ();
 decap_12 FILLER_98_53 ();
 decap_12 FILLER_98_65 ();
 fill_4 FILLER_98_77 ();
 fill_2 FILLER_98_81 ();
 fill_1 FILLER_98_83 ();
 decap_12 FILLER_98_85 ();
 decap_12 FILLER_98_97 ();
 decap_12 FILLER_98_109 ();
 decap_12 FILLER_98_121 ();
 fill_4 FILLER_98_133 ();
 fill_2 FILLER_98_137 ();
 fill_1 FILLER_98_139 ();
 decap_12 FILLER_98_141 ();
 decap_12 FILLER_98_153 ();
 decap_12 FILLER_98_165 ();
 decap_12 FILLER_98_177 ();
 fill_4 FILLER_98_189 ();
 fill_2 FILLER_98_193 ();
 fill_1 FILLER_98_195 ();
 decap_12 FILLER_98_197 ();
 decap_12 FILLER_98_209 ();
 decap_12 FILLER_98_221 ();
 decap_12 FILLER_98_233 ();
 fill_4 FILLER_98_245 ();
 fill_2 FILLER_98_249 ();
 fill_1 FILLER_98_251 ();
 decap_12 FILLER_98_253 ();
 decap_12 FILLER_98_265 ();
 decap_12 FILLER_98_277 ();
 decap_12 FILLER_98_289 ();
 fill_4 FILLER_98_301 ();
 fill_2 FILLER_98_305 ();
 fill_1 FILLER_98_307 ();
 decap_12 FILLER_98_309 ();
 decap_12 FILLER_98_321 ();
 decap_12 FILLER_98_333 ();
 decap_12 FILLER_98_345 ();
 fill_4 FILLER_98_357 ();
 fill_2 FILLER_98_361 ();
 fill_1 FILLER_98_363 ();
 decap_12 FILLER_98_365 ();
 decap_12 FILLER_98_377 ();
 decap_12 FILLER_98_389 ();
 decap_12 FILLER_98_401 ();
 fill_4 FILLER_98_413 ();
 fill_2 FILLER_98_417 ();
 fill_1 FILLER_98_419 ();
 decap_12 FILLER_98_421 ();
 decap_12 FILLER_98_433 ();
 decap_12 FILLER_98_445 ();
 decap_12 FILLER_98_457 ();
 fill_4 FILLER_98_469 ();
 fill_2 FILLER_98_473 ();
 fill_1 FILLER_98_475 ();
 decap_12 FILLER_98_477 ();
 decap_12 FILLER_98_489 ();
 decap_12 FILLER_98_501 ();
 decap_12 FILLER_98_513 ();
 fill_4 FILLER_98_525 ();
 fill_2 FILLER_98_529 ();
 fill_1 FILLER_98_531 ();
 decap_12 FILLER_98_533 ();
 decap_12 FILLER_98_545 ();
 decap_12 FILLER_98_557 ();
 decap_12 FILLER_98_569 ();
 fill_4 FILLER_98_581 ();
 fill_2 FILLER_98_585 ();
 fill_1 FILLER_98_587 ();
 decap_12 FILLER_98_589 ();
 decap_12 FILLER_98_601 ();
 decap_12 FILLER_98_613 ();
 decap_12 FILLER_99_3 ();
 decap_12 FILLER_99_15 ();
 decap_12 FILLER_99_27 ();
 decap_12 FILLER_99_39 ();
 fill_4 FILLER_99_51 ();
 fill_1 FILLER_99_55 ();
 decap_12 FILLER_99_57 ();
 decap_12 FILLER_99_69 ();
 decap_12 FILLER_99_81 ();
 decap_12 FILLER_99_93 ();
 fill_4 FILLER_99_105 ();
 fill_2 FILLER_99_109 ();
 fill_1 FILLER_99_111 ();
 decap_12 FILLER_99_113 ();
 decap_12 FILLER_99_125 ();
 decap_12 FILLER_99_137 ();
 decap_12 FILLER_99_149 ();
 fill_4 FILLER_99_161 ();
 fill_2 FILLER_99_165 ();
 fill_1 FILLER_99_167 ();
 decap_12 FILLER_99_169 ();
 decap_12 FILLER_99_181 ();
 decap_12 FILLER_99_193 ();
 decap_12 FILLER_99_205 ();
 fill_4 FILLER_99_217 ();
 fill_2 FILLER_99_221 ();
 fill_1 FILLER_99_223 ();
 decap_12 FILLER_99_225 ();
 decap_12 FILLER_99_237 ();
 decap_12 FILLER_99_249 ();
 decap_12 FILLER_99_261 ();
 fill_4 FILLER_99_273 ();
 fill_2 FILLER_99_277 ();
 fill_1 FILLER_99_279 ();
 decap_12 FILLER_99_281 ();
 decap_12 FILLER_99_293 ();
 decap_12 FILLER_99_305 ();
 decap_12 FILLER_99_317 ();
 fill_4 FILLER_99_329 ();
 fill_2 FILLER_99_333 ();
 fill_1 FILLER_99_335 ();
 decap_12 FILLER_99_337 ();
 decap_12 FILLER_99_349 ();
 decap_12 FILLER_99_361 ();
 decap_12 FILLER_99_373 ();
 fill_4 FILLER_99_385 ();
 fill_2 FILLER_99_389 ();
 fill_1 FILLER_99_391 ();
 decap_12 FILLER_99_393 ();
 decap_12 FILLER_99_405 ();
 decap_12 FILLER_99_417 ();
 decap_12 FILLER_99_429 ();
 fill_4 FILLER_99_441 ();
 fill_2 FILLER_99_445 ();
 fill_1 FILLER_99_447 ();
 decap_12 FILLER_99_449 ();
 decap_12 FILLER_99_461 ();
 decap_12 FILLER_99_473 ();
 decap_12 FILLER_99_485 ();
 fill_4 FILLER_99_497 ();
 fill_2 FILLER_99_501 ();
 fill_1 FILLER_99_503 ();
 decap_12 FILLER_99_505 ();
 decap_12 FILLER_99_517 ();
 decap_12 FILLER_99_529 ();
 decap_12 FILLER_99_541 ();
 fill_4 FILLER_99_553 ();
 fill_2 FILLER_99_557 ();
 fill_1 FILLER_99_559 ();
 decap_12 FILLER_99_561 ();
 decap_12 FILLER_99_573 ();
 decap_12 FILLER_99_585 ();
 decap_12 FILLER_99_597 ();
 fill_4 FILLER_99_609 ();
 fill_2 FILLER_99_613 ();
 fill_1 FILLER_99_615 ();
 fill_8 FILLER_99_617 ();
 decap_12 FILLER_100_3 ();
 decap_12 FILLER_100_15 ();
 fill_1 FILLER_100_27 ();
 decap_12 FILLER_100_29 ();
 decap_12 FILLER_100_41 ();
 decap_12 FILLER_100_53 ();
 decap_12 FILLER_100_65 ();
 fill_4 FILLER_100_77 ();
 fill_2 FILLER_100_81 ();
 fill_1 FILLER_100_83 ();
 decap_12 FILLER_100_85 ();
 decap_12 FILLER_100_97 ();
 decap_12 FILLER_100_109 ();
 decap_12 FILLER_100_121 ();
 fill_4 FILLER_100_133 ();
 fill_2 FILLER_100_137 ();
 fill_1 FILLER_100_139 ();
 decap_12 FILLER_100_141 ();
 decap_12 FILLER_100_153 ();
 decap_12 FILLER_100_165 ();
 decap_12 FILLER_100_177 ();
 fill_4 FILLER_100_189 ();
 fill_2 FILLER_100_193 ();
 fill_1 FILLER_100_195 ();
 decap_12 FILLER_100_197 ();
 decap_12 FILLER_100_209 ();
 decap_12 FILLER_100_221 ();
 decap_12 FILLER_100_233 ();
 fill_4 FILLER_100_245 ();
 fill_2 FILLER_100_249 ();
 fill_1 FILLER_100_251 ();
 decap_12 FILLER_100_253 ();
 decap_12 FILLER_100_265 ();
 decap_12 FILLER_100_277 ();
 decap_12 FILLER_100_289 ();
 fill_4 FILLER_100_301 ();
 fill_2 FILLER_100_305 ();
 fill_1 FILLER_100_307 ();
 decap_12 FILLER_100_309 ();
 decap_12 FILLER_100_321 ();
 decap_12 FILLER_100_333 ();
 decap_12 FILLER_100_345 ();
 fill_4 FILLER_100_357 ();
 fill_2 FILLER_100_361 ();
 fill_1 FILLER_100_363 ();
 decap_12 FILLER_100_365 ();
 decap_12 FILLER_100_377 ();
 decap_12 FILLER_100_389 ();
 decap_12 FILLER_100_401 ();
 fill_4 FILLER_100_413 ();
 fill_2 FILLER_100_417 ();
 fill_1 FILLER_100_419 ();
 decap_12 FILLER_100_421 ();
 decap_12 FILLER_100_433 ();
 decap_12 FILLER_100_445 ();
 decap_12 FILLER_100_457 ();
 fill_4 FILLER_100_469 ();
 fill_2 FILLER_100_473 ();
 fill_1 FILLER_100_475 ();
 decap_12 FILLER_100_477 ();
 decap_12 FILLER_100_489 ();
 decap_12 FILLER_100_501 ();
 decap_12 FILLER_100_513 ();
 fill_4 FILLER_100_525 ();
 fill_2 FILLER_100_529 ();
 fill_1 FILLER_100_531 ();
 decap_12 FILLER_100_533 ();
 decap_12 FILLER_100_545 ();
 decap_12 FILLER_100_557 ();
 decap_12 FILLER_100_569 ();
 fill_4 FILLER_100_581 ();
 fill_2 FILLER_100_585 ();
 fill_1 FILLER_100_587 ();
 decap_12 FILLER_100_589 ();
 decap_12 FILLER_100_601 ();
 decap_12 FILLER_100_613 ();
 decap_12 FILLER_101_3 ();
 decap_12 FILLER_101_15 ();
 fill_1 FILLER_101_27 ();
 decap_12 FILLER_101_29 ();
 decap_12 FILLER_101_41 ();
 fill_2 FILLER_101_53 ();
 fill_1 FILLER_101_55 ();
 decap_12 FILLER_101_57 ();
 decap_12 FILLER_101_69 ();
 fill_2 FILLER_101_81 ();
 fill_1 FILLER_101_83 ();
 decap_12 FILLER_101_85 ();
 decap_12 FILLER_101_97 ();
 fill_2 FILLER_101_109 ();
 fill_1 FILLER_101_111 ();
 decap_12 FILLER_101_113 ();
 decap_12 FILLER_101_125 ();
 fill_2 FILLER_101_137 ();
 fill_1 FILLER_101_139 ();
 decap_12 FILLER_101_141 ();
 decap_12 FILLER_101_153 ();
 fill_2 FILLER_101_165 ();
 fill_1 FILLER_101_167 ();
 decap_12 FILLER_101_169 ();
 decap_12 FILLER_101_181 ();
 fill_2 FILLER_101_193 ();
 fill_1 FILLER_101_195 ();
 decap_12 FILLER_101_197 ();
 decap_12 FILLER_101_209 ();
 fill_2 FILLER_101_221 ();
 fill_1 FILLER_101_223 ();
 decap_12 FILLER_101_225 ();
 decap_12 FILLER_101_237 ();
 fill_2 FILLER_101_249 ();
 fill_1 FILLER_101_251 ();
 decap_12 FILLER_101_253 ();
 decap_12 FILLER_101_265 ();
 fill_2 FILLER_101_277 ();
 fill_1 FILLER_101_279 ();
 decap_12 FILLER_101_281 ();
 decap_12 FILLER_101_293 ();
 fill_2 FILLER_101_305 ();
 fill_1 FILLER_101_307 ();
 decap_12 FILLER_101_309 ();
 decap_12 FILLER_101_321 ();
 fill_2 FILLER_101_333 ();
 fill_1 FILLER_101_335 ();
 decap_12 FILLER_101_337 ();
 decap_12 FILLER_101_349 ();
 fill_2 FILLER_101_361 ();
 fill_1 FILLER_101_363 ();
 decap_12 FILLER_101_365 ();
 decap_12 FILLER_101_377 ();
 fill_2 FILLER_101_389 ();
 fill_1 FILLER_101_391 ();
 decap_12 FILLER_101_393 ();
 decap_12 FILLER_101_405 ();
 fill_2 FILLER_101_417 ();
 fill_1 FILLER_101_419 ();
 decap_12 FILLER_101_421 ();
 decap_12 FILLER_101_433 ();
 fill_2 FILLER_101_445 ();
 fill_1 FILLER_101_447 ();
 decap_12 FILLER_101_449 ();
 decap_12 FILLER_101_461 ();
 fill_2 FILLER_101_473 ();
 fill_1 FILLER_101_475 ();
 decap_12 FILLER_101_477 ();
 decap_12 FILLER_101_489 ();
 fill_2 FILLER_101_501 ();
 fill_1 FILLER_101_503 ();
 decap_12 FILLER_101_505 ();
 decap_12 FILLER_101_517 ();
 fill_2 FILLER_101_529 ();
 fill_1 FILLER_101_531 ();
 decap_12 FILLER_101_533 ();
 decap_12 FILLER_101_545 ();
 fill_2 FILLER_101_557 ();
 fill_1 FILLER_101_559 ();
 decap_12 FILLER_101_561 ();
 decap_12 FILLER_101_573 ();
 fill_2 FILLER_101_585 ();
 fill_1 FILLER_101_587 ();
 decap_12 FILLER_101_589 ();
 decap_12 FILLER_101_601 ();
 fill_2 FILLER_101_613 ();
 fill_1 FILLER_101_615 ();
 fill_8 FILLER_101_617 ();

endmodule
