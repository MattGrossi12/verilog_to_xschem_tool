module digitop_pav2_mpw03 (
    input clk_i,
    input demod_i,
    input rnclk_i,
    input [63:0] rr_data_i,
    input rst_b_i,
    input se_i,
    input sel_nvm_i,
    input tclk_i,
    input ti_i,
    output amux_en_o,
    output amux_ib_sel_o,
    output amux_vcc_sel_o,
    output amux_vdd_sel_o,
    output amux_vref_sel_o,
    output [2:0] clk_trim_o,
    output demod_en_o,
    output mod_o,
    output rnclk_en_o,
    output [2:0] rnclk_trim_o,
    output [3:0] rr_bank_sel_o,
    output [15:0] rr_bl_o,
    output rr_erase_o,
    output rr_form_en_o,
    output rr_prog_o,
    output rr_read_o,
    output [31:0] rr_wl_o,
    output to_dig_en_b_o,
    output to_o
);

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire \digitop_pav2.acc_activate ;
 wire \digitop_pav2.access_inst.acc_wcknzero_o ;
 wire \digitop_pav2.access_inst.access_check0.act_lock_st ;
 wire \digitop_pav2.access_inst.access_check0.clk_i ;
 wire \digitop_pav2.access_inst.access_check0.ctrl_wcknzero_ck ;
 wire \digitop_pav2.access_inst.access_check0.error_word_cnt_ptr ;
 wire \digitop_pav2.access_inst.access_check0.error_wordcnt_i ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[0] ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[10] ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[11] ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[13] ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[1] ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[2] ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[3] ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[4] ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[5] ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[6] ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[7] ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[8] ;
 wire \digitop_pav2.access_inst.access_check0.fg_i[9] ;
 wire \digitop_pav2.access_inst.access_check0.g_activate_i ;
 wire \digitop_pav2.access_inst.access_check0.g_propwrite_i ;
 wire \digitop_pav2.access_inst.access_check0.g_read_i ;
 wire \digitop_pav2.access_inst.access_check0.g_write_i ;
 wire \digitop_pav2.access_inst.access_check0.lock_error_o ;
 wire \digitop_pav2.access_inst.access_check0.mem_sign_check_i ;
 wire \digitop_pav2.access_inst.access_check0.mem_sign_check_sync_o ;
 wire \digitop_pav2.access_inst.access_check0.pc_invalid_o ;
 wire \digitop_pav2.access_inst.access_check0.pc_lock_check_i ;
 wire \digitop_pav2.access_inst.access_check0.pc_lock_check_sync_o ;
 wire \digitop_pav2.access_inst.access_check0.permalock_tid_i ;
 wire \digitop_pav2.access_inst.access_check0.proc_finish1_i ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[0] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[10] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[11] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[12] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[13] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[14] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[15] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[1] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[2] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[3] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[4] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[5] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[6] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[7] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[8] ;
 wire \digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[9] ;
 wire \digitop_pav2.access_inst.access_check0.wcnt_check_one ;
 wire \digitop_pav2.access_inst.access_check0.wcnt_check_zero ;
 wire \digitop_pav2.access_inst.access_check0.wordcnt_i[0] ;
 wire \digitop_pav2.access_inst.access_check0.wordcnt_i[1] ;
 wire \digitop_pav2.access_inst.access_check0.wordcnt_i[2] ;
 wire \digitop_pav2.access_inst.access_check0.wordcnt_i[3] ;
 wire \digitop_pav2.access_inst.access_check0.wordcnt_i[4] ;
 wire \digitop_pav2.access_inst.access_check0.wordcnt_i[5] ;
 wire \digitop_pav2.access_inst.access_check0.wordcnt_i[6] ;
 wire \digitop_pav2.access_inst.access_check0.wordptr_i[0] ;
 wire \digitop_pav2.access_inst.access_check0.wordptr_i[1] ;
 wire \digitop_pav2.access_inst.access_check0.wordptr_i[2] ;
 wire \digitop_pav2.access_inst.access_check0.wordptr_i[3] ;
 wire \digitop_pav2.access_inst.access_check0.wordptr_i[4] ;
 wire \digitop_pav2.access_inst.access_check0.wordptr_i[5] ;
 wire \digitop_pav2.access_inst.access_check0.wordptr_i[6] ;
 wire \digitop_pav2.access_inst.access_check0.wr_check_sync_o ;
 wire \digitop_pav2.access_inst.access_check0.wr_key_ck_i ;
 wire \digitop_pav2.access_inst.access_check0.wr_lock_ck_i ;
 wire \digitop_pav2.access_inst.access_check0.write_check_i ;
 wire \digitop_pav2.access_inst.access_check0.write_error_reg ;
 wire \digitop_pav2.access_inst.access_ctrl0.crc_en_o ;
 wire \digitop_pav2.access_inst.access_ctrl0.crc_init_i ;
 wire \digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt ;
 wire \digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt_ok ;
 wire \digitop_pav2.access_inst.access_ctrl0.dt_acc_done ;
 wire \digitop_pav2.access_inst.access_ctrl0.dt_acc_done_o ;
 wire \digitop_pav2.access_inst.access_ctrl0.f_access_i ;
 wire \digitop_pav2.access_inst.access_ctrl0.ld_dt_env_finish_i ;
 wire \digitop_pav2.access_inst.access_ctrl0.ld_dt_stb ;
 wire \digitop_pav2.access_inst.access_ctrl0.ld_key_env_finish_i ;
 wire \digitop_pav2.access_inst.access_ctrl0.nvm_busy_i ;
 wire \digitop_pav2.access_inst.access_ctrl0.prev_busy ;
 wire \digitop_pav2.access_inst.access_ctrl0.proc_finish0_i ;
 wire \digitop_pav2.access_inst.access_ctrl0.proc_rd_finish_i ;
 wire \digitop_pav2.access_inst.access_ctrl0.replay_nok ;
 wire \digitop_pav2.access_inst.access_ctrl0.replay_ok ;
 wire \digitop_pav2.access_inst.access_ctrl0.rx_par0_i ;
 wire \digitop_pav2.access_inst.access_ctrl0.rx_par1_i ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[0] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[10] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[11] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[13] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[14] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[15] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[17] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[18] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[19] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[1] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[20] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[22] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[23] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[24] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[25] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[2] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[5] ;
 wire \digitop_pav2.access_inst.access_ctrl0.state[9] ;
 wire \digitop_pav2.access_inst.access_ctrl0.tx_bit_i ;
 wire \digitop_pav2.access_inst.access_ctrl0.tx_dt_finish_i ;
 wire \digitop_pav2.access_inst.access_ctrl0.tx_proc_rd_stb_i ;
 wire \digitop_pav2.access_inst.access_ctrl0.wr_key_finish_i ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[0] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[10] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[11] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[12] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[13] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[14] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[15] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[1] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[2] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[3] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[4] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[5] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[6] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[7] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[8] ;
 wire \digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[9] ;
 wire \digitop_pav2.access_inst.access_proc0.ctrl_rd_bus ;
 wire \digitop_pav2.access_inst.access_proc0.ctrl_rd_bus_res ;
 wire \digitop_pav2.access_inst.access_proc0.nvm_acc_addr[0] ;
 wire \digitop_pav2.access_inst.access_proc0.nvm_acc_addr[1] ;
 wire \digitop_pav2.access_inst.access_proc0.nvm_acc_addr[2] ;
 wire \digitop_pav2.access_inst.access_proc0.nvm_acc_addr[3] ;
 wire \digitop_pav2.access_inst.access_proc0.nvm_acc_addr[4] ;
 wire \digitop_pav2.access_inst.access_proc0.nvm_acc_addr[5] ;
 wire \digitop_pav2.access_inst.access_proc0.nvm_acc_addr[6] ;
 wire \digitop_pav2.access_inst.access_proc0.nvm_acc_addr[7] ;
 wire \digitop_pav2.access_inst.access_proc0.nvm_acc_addr[8] ;
 wire \digitop_pav2.access_inst.access_proc0.proc_crc_check[0] ;
 wire \digitop_pav2.access_inst.access_proc0.proc_crc_check[1] ;
 wire \digitop_pav2.access_inst.access_proc0.proc_crc_check[2] ;
 wire \digitop_pav2.access_inst.access_proc0.proc_crc_check[3] ;
 wire \digitop_pav2.access_inst.access_proc0.proc_crc_check[4] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[0] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[10] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[11] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[12] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[13] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[14] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[15] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[1] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[2] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[3] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[4] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[5] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[6] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[7] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[8] ;
 wire \digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[9] ;
 wire \digitop_pav2.access_inst.access_transceiver0.ctrl_circ_buf ;
 wire \digitop_pav2.access_inst.access_transceiver0.dt_ptr[0] ;
 wire \digitop_pav2.access_inst.access_transceiver0.dt_ptr[1] ;
 wire \digitop_pav2.access_inst.access_transceiver0.dt_ptr[2] ;
 wire \digitop_pav2.access_inst.access_transceiver0.dt_ptr[3] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[0] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[10] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[11] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[12] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[13] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[14] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[15] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[1] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[2] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[3] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[4] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[5] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[6] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[7] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[8] ;
 wire \digitop_pav2.access_inst.access_transceiver0.handle_i[9] ;
 wire \digitop_pav2.access_inst.access_transceiver0.rx_par_buf[14] ;
 wire \digitop_pav2.access_inst.access_transceiver0.rx_par_buf[15] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[0] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[10] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[11] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[12] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[13] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[14] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[15] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[1] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[2] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[3] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[4] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[5] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[6] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[7] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[8] ;
 wire \digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[9] ;
 wire \digitop_pav2.access_inst.access_transceiver0.wcnt_stb_valid ;
 wire \digitop_pav2.ack_inst.buffer_ff[0] ;
 wire \digitop_pav2.ack_inst.buffer_ff[10] ;
 wire \digitop_pav2.ack_inst.buffer_ff[11] ;
 wire \digitop_pav2.ack_inst.buffer_ff[12] ;
 wire \digitop_pav2.ack_inst.buffer_ff[13] ;
 wire \digitop_pav2.ack_inst.buffer_ff[14] ;
 wire \digitop_pav2.ack_inst.buffer_ff[15] ;
 wire \digitop_pav2.ack_inst.buffer_ff[1] ;
 wire \digitop_pav2.ack_inst.buffer_ff[2] ;
 wire \digitop_pav2.ack_inst.buffer_ff[3] ;
 wire \digitop_pav2.ack_inst.buffer_ff[4] ;
 wire \digitop_pav2.ack_inst.buffer_ff[5] ;
 wire \digitop_pav2.ack_inst.buffer_ff[6] ;
 wire \digitop_pav2.ack_inst.buffer_ff[7] ;
 wire \digitop_pav2.ack_inst.buffer_ff[8] ;
 wire \digitop_pav2.ack_inst.buffer_ff[9] ;
 wire \digitop_pav2.ack_inst.clk_i ;
 wire \digitop_pav2.ack_inst.cnt_ff[0] ;
 wire \digitop_pav2.ack_inst.cnt_ff[1] ;
 wire \digitop_pav2.ack_inst.cnt_ff[2] ;
 wire \digitop_pav2.ack_inst.cnt_ff[3] ;
 wire \digitop_pav2.ack_inst.g_ack_i ;
 wire \digitop_pav2.ack_inst.nvm_ack_rd_stb_o ;
 wire \digitop_pav2.ack_inst.rcnt_ff[0] ;
 wire \digitop_pav2.ack_inst.rcnt_ff[1] ;
 wire \digitop_pav2.ack_inst.state_ff[0] ;
 wire \digitop_pav2.ack_inst.state_ff[1] ;
 wire \digitop_pav2.ack_inst.state_ff[2] ;
 wire \digitop_pav2.aes128_inst.aes128_counter.clk_i ;
 wire \digitop_pav2.aes128_inst.aes128_counter.cnt_fin_2b_o ;
 wire \digitop_pav2.aes128_inst.aes128_counter.cnt_fin_3b_o ;
 wire \digitop_pav2.aes128_inst.aes128_counter.cnt_fin_key_o ;
 wire \digitop_pav2.aes128_inst.aes128_counter.cnt_rnd_en_o ;
 wire \digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[0] ;
 wire \digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[1] ;
 wire \digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[2] ;
 wire \digitop_pav2.aes128_inst.aes128_counter.rst_b_i ;
 wire \digitop_pav2.aes128_inst.aes128_regs.aes_exe_o ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key0_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key1_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key2_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key3_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key4_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key5_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key6_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.key7_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.rcon_i[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.rcon_i[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.rcon_i[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.rcon_i[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.rcon_i[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.rcon_i[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.rcon_i[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.rcon_i[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state0_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state1_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state2_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state3_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state4_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state5_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state6_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[10] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[11] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[12] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[13] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[14] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[15] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[8] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state7_r[9] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state_areg_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state_areg_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state_areg_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state_areg_r[3] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state_areg_r[4] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state_areg_r[5] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state_areg_r[6] ;
 wire \digitop_pav2.aes128_inst.aes128_regs.state_areg_r[7] ;
 wire \digitop_pav2.aes128_inst.aes128_round.round_cnt_r[0] ;
 wire \digitop_pav2.aes128_inst.aes128_round.round_cnt_r[1] ;
 wire \digitop_pav2.aes128_inst.aes128_round.round_cnt_r[2] ;
 wire \digitop_pav2.aes128_inst.aes128_round.round_cnt_r[3] ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_0.A ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_0.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_1.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_2.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_3.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_4.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_5.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_6.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_7.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_8.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_9.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_0.A ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_0.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_1.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_2.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_3.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_4.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_5.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_6.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_7.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_8.Y ;
 wire \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_9.Y ;
 wire \digitop_pav2.boot_inst.boot_ctrl0.act_state_i ;
 wire \digitop_pav2.boot_inst.boot_ctrl0.clk_i ;
 wire \digitop_pav2.boot_inst.boot_ctrl0.ctrl_crc_en ;
 wire \digitop_pav2.boot_inst.boot_ctrl0.ctrl_replay_o ;
 wire \digitop_pav2.boot_inst.boot_ctrl0.prev_busy ;
 wire \digitop_pav2.boot_inst.boot_ctrl0.proc_boot_end_i ;
 wire \digitop_pav2.boot_inst.boot_ctrl0.proc_crc_end_i ;
 wire \digitop_pav2.boot_inst.boot_ctrl0.replay ;
 wire \digitop_pav2.boot_inst.boot_ctrl0.state[0] ;
 wire \digitop_pav2.boot_inst.boot_ctrl0.state[2] ;
 wire \digitop_pav2.boot_inst.boot_ctrl0.state[3] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[0] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[10] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[11] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[12] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[13] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[14] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[15] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[1] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[2] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[3] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[4] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[5] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[6] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[7] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[8] ;
 wire \digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[9] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_boot_sync ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_fg[12] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[0] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[10] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[11] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[12] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[13] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[14] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[15] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[16] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[17] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[18] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[19] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[1] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[20] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[21] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[22] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[23] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[24] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[25] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[26] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[27] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[28] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[29] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[2] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[30] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[31] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[3] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[4] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[5] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[6] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[7] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[8] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_mask[9] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_stage[0] ;
 wire \digitop_pav2.boot_inst.boot_proc0.proc_stage[1] ;
 wire \digitop_pav2.boot_inst.r_boot_ff ;
 wire \digitop_pav2.cal_inst.calx_clk_o ;
 wire \digitop_pav2.cal_inst.calx_mux.dtest_trim_0_i ;
 wire \digitop_pav2.cal_inst.calx_mux.dtest_trim_1_i ;
 wire \digitop_pav2.cal_inst.calx_mux.dtest_trim_2_i ;
 wire \digitop_pav2.cal_inst.calx_mux.en_calx_test_i ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.aux_clk ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.auxclk_after_buf ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.ck_in ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.ck_out ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.enable ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.w_nor ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.w_not ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk2 ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk2_after_buf ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk4 ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk_dftmux.dft_rp_and ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.end_stab_clk_i ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.ref_pulse_sync_o ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.rp_ff[0] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_clk.stab_clk_dis ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.calx_end_o ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.en_pctr ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_end ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_end_stab_clk ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_rd_stb ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_state[0] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_state[1] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_state[2] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_state[3] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_wr_stb ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.nvm_calx_rd_stb_o ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.nvm_calx_wr_stb_o ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[0] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[1] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[2] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[3] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[4] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[5] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[6] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[7] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[8] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[9] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[0] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[1] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[2] ;
 wire \digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[3] ;
 wire \digitop_pav2.clkx_cp_clk ;
 wire \digitop_pav2.clkx_fm0x_clk ;
 wire \digitop_pav2.clkx_invent_clk ;
 wire \digitop_pav2.clkx_irreg_clk ;
 wire \digitop_pav2.clkx_mem_top_clk ;
 wire \digitop_pav2.clkx_past_irreg_clk ;
 wire \digitop_pav2.clkx_piex_clk ;
 wire \digitop_pav2.clkx_rngx_clk ;
 wire \digitop_pav2.clkx_rngx_fast_clk ;
 wire \digitop_pav2.clkx_sec_clk ;
 wire \digitop_pav2.crc_eval ;
 wire \digitop_pav2.crc_inst.count[0] ;
 wire \digitop_pav2.crc_inst.count[1] ;
 wire \digitop_pav2.crc_inst.count[2] ;
 wire \digitop_pav2.crc_inst.count[3] ;
 wire \digitop_pav2.crc_inst.crc16_q[0] ;
 wire \digitop_pav2.crc_inst.crc16_q[10] ;
 wire \digitop_pav2.crc_inst.crc16_q[11] ;
 wire \digitop_pav2.crc_inst.crc16_q[12] ;
 wire \digitop_pav2.crc_inst.crc16_q[13] ;
 wire \digitop_pav2.crc_inst.crc16_q[14] ;
 wire \digitop_pav2.crc_inst.crc16_q[15] ;
 wire \digitop_pav2.crc_inst.crc16_q[1] ;
 wire \digitop_pav2.crc_inst.crc16_q[2] ;
 wire \digitop_pav2.crc_inst.crc16_q[3] ;
 wire \digitop_pav2.crc_inst.crc16_q[4] ;
 wire \digitop_pav2.crc_inst.crc16_q[5] ;
 wire \digitop_pav2.crc_inst.crc16_q[6] ;
 wire \digitop_pav2.crc_inst.crc16_q[7] ;
 wire \digitop_pav2.crc_inst.crc16_q[8] ;
 wire \digitop_pav2.crc_inst.crc16_q[9] ;
 wire \digitop_pav2.crc_inst.crc5_q[0] ;
 wire \digitop_pav2.crc_inst.crc5_q[1] ;
 wire \digitop_pav2.crc_inst.crc5_q[2] ;
 wire \digitop_pav2.crc_inst.crc5_q[3] ;
 wire \digitop_pav2.crc_inst.crc5_q[4] ;
 wire \digitop_pav2.crc_inst.dt_rx_en_i ;
 wire \digitop_pav2.crc_inst.dt_rx_i ;
 wire \digitop_pav2.crc_inst.dt_tx_en_aux ;
 wire \digitop_pav2.crc_inst.mctrl_data_en_ff ;
 wire \digitop_pav2.crc_inst.mctrl_data_end_ff ;
 wire \digitop_pav2.crc_inst.pie_data_en_ff ;
 wire \digitop_pav2.dr ;
 wire \digitop_pav2.fg_tc ;
 wire \digitop_pav2.fm0miller_inst.ctrl[0] ;
 wire \digitop_pav2.fm0miller_inst.ctrl[1] ;
 wire \digitop_pav2.fm0miller_inst.ctrl[2] ;
 wire \digitop_pav2.fm0miller_inst.dt_tx_st_o ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[0] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[1] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[2] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[3] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[4] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[0] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[1] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[2] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[3] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[4] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[5] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[6] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[0] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[1] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[2] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[3] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[4] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[5] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[6] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.en_i ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[0] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[1] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[2] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.mod_en ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.n_data_valid ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.n_dt_tx_st ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.n_gand ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.n_gor ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.state[0] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.state[1] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_ctrl.state[2] ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.gand ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.gand_delay ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[0].fm0miller_pav2_gand_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[0].fm0miller_pav2_gor_dly.A ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[0].fm0miller_pav2_gor_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[1].fm0miller_pav2_gand_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[1].fm0miller_pav2_gor_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[2].fm0miller_pav2_gand_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[2].fm0miller_pav2_gor_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[3].fm0miller_pav2_gand_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[3].fm0miller_pav2_gor_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[4].fm0miller_pav2_gand_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[4].fm0miller_pav2_gor_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[5].fm0miller_pav2_gand_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[5].fm0miller_pav2_gor_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[6].fm0miller_pav2_gand_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[6].fm0miller_pav2_gor_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[7].fm0miller_pav2_gand_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[7].fm0miller_pav2_gor_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[8].fm0miller_pav2_gand_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[8].fm0miller_pav2_gor_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[9].fm0miller_pav2_gor_dly.Y ;
 wire \digitop_pav2.fm0miller_inst.fm0x_mask.tx_raw_i ;
 wire net1610;
 wire net1617;
 wire \digitop_pav2.fm0miller_inst.fm0x_tx.data_fm0x_clk_is_data_after_buf ;
 wire \digitop_pav2.fm0miller_inst.fm0x_tx.data_fm0x_clk_is_data_after_buf_b ;
 wire \digitop_pav2.fm0miller_inst.fm0x_tx.w_fmdata_mux_0 ;
 wire \digitop_pav2.fm0miller_inst.fm0x_tx.w_fmdata_mux_1 ;
 wire \digitop_pav2.fm0x_clk_for_proc_ctrl ;
 wire \digitop_pav2.func_clk ;
 wire \digitop_pav2.func_clk_pre ;
 wire \digitop_pav2.func_reg_wr_en ;
 wire \digitop_pav2.func_rnclk_en ;
 wire \digitop_pav2.func_rng_data[0] ;
 wire \digitop_pav2.func_rng_data[10] ;
 wire \digitop_pav2.func_rng_data[11] ;
 wire \digitop_pav2.func_rng_data[12] ;
 wire \digitop_pav2.func_rng_data[13] ;
 wire \digitop_pav2.func_rng_data[14] ;
 wire \digitop_pav2.func_rng_data[15] ;
 wire \digitop_pav2.func_rng_data[1] ;
 wire \digitop_pav2.func_rng_data[2] ;
 wire \digitop_pav2.func_rng_data[3] ;
 wire \digitop_pav2.func_rng_data[4] ;
 wire \digitop_pav2.func_rng_data[5] ;
 wire \digitop_pav2.func_rng_data[6] ;
 wire \digitop_pav2.func_rng_data[7] ;
 wire \digitop_pav2.func_rng_data[8] ;
 wire \digitop_pav2.func_rng_data[9] ;
 wire \digitop_pav2.func_rr_erase ;
 wire \digitop_pav2.func_rr_prog ;
 wire \digitop_pav2.func_rr_read ;
 wire \digitop_pav2.g_auth_obu ;
 wire \digitop_pav2.g_query ;
 wire \digitop_pav2.g_queryadj ;
 wire \digitop_pav2.g_queryrep ;
 wire \digitop_pav2.g_reqrn ;
 wire \digitop_pav2.g_select ;
 wire \digitop_pav2.glue_inst.mbus_rd_en_o ;
 wire \digitop_pav2.glue_inst.mbus_wr_en_o ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[1] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[2] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[3] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[4] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[5] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[6] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[7] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[0] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[1] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[2] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[3] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[4] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[5] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[6] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[7] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[0] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[1] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[2] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[3] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[4] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[5] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[6] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[7] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[0] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[1] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[2] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[3] ;
 wire \digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[4] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.flags_en_o ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[0] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[1] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.q[0] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.q[1] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.q[2] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.q[3] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.query_inversion ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.r_invent2_o ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.r_invent3_o ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.s0_i ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.s1_i ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.s2_i ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.s2_r_ff_i ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.s2_s_ff_i ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.s3_r_ff_i ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.s3_s_ff_i ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.sl_i ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[0] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[10] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[11] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[12] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[13] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[14] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[1] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[2] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[3] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[4] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[5] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[6] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[7] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[8] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[9] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.state[0] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.state[11] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.state[13] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.state[1] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.state[2] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.state[3] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.state[4] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.state[5] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.state[6] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.state[7] ;
 wire \digitop_pav2.invent_inst.invent_qqqr_pav2.state[9] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.bitptr[0] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.bitptr[1] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.bitptr[2] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.bitptr[3] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.bitptr[4] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.bitptr[5] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.bitptr[6] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.bitptr[7] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.bitptr[8] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[0] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[10] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[11] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[12] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[13] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[14] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[15] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[1] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[2] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[3] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[4] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[5] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[6] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[7] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[8] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf1[9] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[0] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[10] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[11] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[12] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[13] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[14] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[15] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[1] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[2] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[3] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[4] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[5] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[6] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[7] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[8] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.buf2[9] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.mask_mismatch_ff ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.r_invent2_o ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.r_invent3_o ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.select_valid_o ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.state[0] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.state[10] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.state[11] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.state[12] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.state[1] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.state[2] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.state[4] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.state[5] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.state[6] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.state[7] ;
 wire \digitop_pav2.invent_inst.invent_sel_pav2.state[9] ;
 wire \digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[0] ;
 wire \digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[1] ;
 wire \digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[2] ;
 wire \digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[3] ;
 wire \digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[4] ;
 wire \digitop_pav2.invent_inst.s1_i ;
 wire \digitop_pav2.invent_inst.s1_r_o ;
 wire \digitop_pav2.invent_inst.s1_s_o ;
 wire \digitop_pav2.invent_inst.s2_r_o ;
 wire \digitop_pav2.invent_inst.s2_s_o ;
 wire \digitop_pav2.invent_inst.s3_r_o ;
 wire \digitop_pav2.invent_inst.s3_s_o ;
 wire \digitop_pav2.invent_inst.sl_r_ff ;
 wire \digitop_pav2.invent_inst.sl_r_o ;
 wire \digitop_pav2.invent_inst.sl_s_ff ;
 wire \digitop_pav2.invent_inst.sl_s_o ;
 wire \digitop_pav2.memctrl_inst.addr_to_reram[0] ;
 wire \digitop_pav2.memctrl_inst.addr_to_reram[1] ;
 wire \digitop_pav2.memctrl_inst.addr_to_reram[2] ;
 wire \digitop_pav2.memctrl_inst.addr_to_reram[3] ;
 wire \digitop_pav2.memctrl_inst.addr_to_reram[4] ;
 wire \digitop_pav2.memctrl_inst.bit_addr[0] ;
 wire \digitop_pav2.memctrl_inst.bit_addr[1] ;
 wire \digitop_pav2.memctrl_inst.bit_addr[2] ;
 wire \digitop_pav2.memctrl_inst.bit_addr[3] ;
 wire \digitop_pav2.memctrl_inst.bit_addr_allow ;
 wire \digitop_pav2.memctrl_inst.busy_ff ;
 wire \digitop_pav2.memctrl_inst.ctr[0] ;
 wire \digitop_pav2.memctrl_inst.ctr[1] ;
 wire \digitop_pav2.memctrl_inst.ctr[2] ;
 wire \digitop_pav2.memctrl_inst.ctr[3] ;
 wire \digitop_pav2.memctrl_inst.ctr[4] ;
 wire \digitop_pav2.memctrl_inst.ctr[5] ;
 wire \digitop_pav2.memctrl_inst.ctr[6] ;
 wire \digitop_pav2.memctrl_inst.ctr[7] ;
 wire \digitop_pav2.memctrl_inst.extra_dt_i[12] ;
 wire \digitop_pav2.memctrl_inst.extra_dt_i[13] ;
 wire \digitop_pav2.memctrl_inst.extra_dt_i[14] ;
 wire \digitop_pav2.memctrl_inst.extra_dt_i[15] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[0] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[10] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[11] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[12] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[13] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[14] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[15] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[1] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[2] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[3] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[4] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[5] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[6] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[7] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[8] ;
 wire \digitop_pav2.memctrl_inst.flops_0x081[9] ;
 wire \digitop_pav2.memctrl_inst.n_bit_addr_allow ;
 wire \digitop_pav2.memctrl_inst.n_erase ;
 wire \digitop_pav2.memctrl_inst.n_prog ;
 wire \digitop_pav2.memctrl_inst.n_read ;
 wire \digitop_pav2.memctrl_inst.n_state[2] ;
 wire \digitop_pav2.memctrl_inst.nvm_rd_en_i ;
 wire \digitop_pav2.memctrl_inst.nvm_wr_en_i ;
 wire \digitop_pav2.memctrl_inst.reg_wr_ok_ff ;
 wire \digitop_pav2.memctrl_inst.reg_wr_ok_ff2 ;
 wire \digitop_pav2.memctrl_inst.state[0] ;
 wire \digitop_pav2.memctrl_inst.state[1] ;
 wire \digitop_pav2.memctrl_inst.state[2] ;
 wire \digitop_pav2.memctrl_inst.state[3] ;
 wire \digitop_pav2.memctrl_inst.state[4] ;
 wire \digitop_pav2.pass_t2 ;
 wire \digitop_pav2.pie_inst.ctr.en_ctr_after_buf ;
 wire \digitop_pav2.pie_inst.ctr.en_ctr_i ;
 wire \digitop_pav2.pie_inst.ctr.ovf_b ;
 wire \digitop_pav2.pie_inst.delend_o ;
 wire \digitop_pav2.pie_inst.en_ctr ;
 wire \digitop_pav2.pie_inst.en_ctr_fix ;
 wire \digitop_pav2.pie_inst.fsm.clk_i ;
 wire \digitop_pav2.pie_inst.fsm.comp_delimiter_ff ;
 wire \digitop_pav2.pie_inst.fsm.comp_delimiter_ff2 ;
 wire \digitop_pav2.pie_inst.fsm.comp_tari_ff ;
 wire \digitop_pav2.pie_inst.fsm.dif_pos_fix[0] ;
 wire \digitop_pav2.pie_inst.fsm.dif_pos_fix[1] ;
 wire \digitop_pav2.pie_inst.fsm.dif_pos_fix[2] ;
 wire \digitop_pav2.pie_inst.fsm.dif_pos_fix[3] ;
 wire \digitop_pav2.pie_inst.fsm.dif_pos_fix[4] ;
 wire \digitop_pav2.pie_inst.fsm.dif_pos_fix[5] ;
 wire \digitop_pav2.pie_inst.fsm.dif_pos_fix[6] ;
 wire \digitop_pav2.pie_inst.fsm.dif_pos_fix[7] ;
 wire \digitop_pav2.pie_inst.fsm.dif_pos_fix[8] ;
 wire \digitop_pav2.pie_inst.fsm.dif_pos_fix[9] ;
 wire \digitop_pav2.pie_inst.fsm.n_data_en ;
 wire \digitop_pav2.pie_inst.fsm.neg_i[1] ;
 wire \digitop_pav2.pie_inst.fsm.neg_i[2] ;
 wire \digitop_pav2.pie_inst.fsm.neg_i[3] ;
 wire \digitop_pav2.pie_inst.fsm.neg_i[4] ;
 wire \digitop_pav2.pie_inst.fsm.neg_i[5] ;
 wire \digitop_pav2.pie_inst.fsm.neg_i[6] ;
 wire \digitop_pav2.pie_inst.fsm.neg_i[7] ;
 wire \digitop_pav2.pie_inst.fsm.neg_i[8] ;
 wire \digitop_pav2.pie_inst.fsm.neg_i[9] ;
 wire \digitop_pav2.pie_inst.fsm.past_clk_i ;
 wire \digitop_pav2.pie_inst.fsm.past_ctr[1] ;
 wire \digitop_pav2.pie_inst.fsm.past_ctr[2] ;
 wire \digitop_pav2.pie_inst.fsm.past_ctr[3] ;
 wire \digitop_pav2.pie_inst.fsm.past_ctr[4] ;
 wire \digitop_pav2.pie_inst.fsm.past_ctr[5] ;
 wire \digitop_pav2.pie_inst.fsm.past_ctr[6] ;
 wire \digitop_pav2.pie_inst.fsm.past_ctr[7] ;
 wire \digitop_pav2.pie_inst.fsm.past_ctr[8] ;
 wire \digitop_pav2.pie_inst.fsm.past_ctr[9] ;
 wire \digitop_pav2.pie_inst.fsm.past_ovf_b ;
 wire \digitop_pav2.pie_inst.fsm.pivot[0] ;
 wire \digitop_pav2.pie_inst.fsm.pivot[1] ;
 wire \digitop_pav2.pie_inst.fsm.pivot[2] ;
 wire \digitop_pav2.pie_inst.fsm.pivot[3] ;
 wire \digitop_pav2.pie_inst.fsm.pivot[4] ;
 wire \digitop_pav2.pie_inst.fsm.pivot[5] ;
 wire \digitop_pav2.pie_inst.fsm.pivot[6] ;
 wire \digitop_pav2.pie_inst.fsm.pivot[7] ;
 wire \digitop_pav2.pie_inst.fsm.pivot[8] ;
 wire \digitop_pav2.pie_inst.fsm.state[0] ;
 wire \digitop_pav2.pie_inst.fsm.state[1] ;
 wire \digitop_pav2.pie_inst.fsm.temptari[0] ;
 wire \digitop_pav2.pie_inst.fsm.temptari[1] ;
 wire \digitop_pav2.pie_inst.fsm.temptari[2] ;
 wire \digitop_pav2.pie_inst.fsm.temptari[3] ;
 wire \digitop_pav2.pie_inst.fsm.temptari[4] ;
 wire \digitop_pav2.pie_inst.fsm.temptari[5] ;
 wire \digitop_pav2.pie_inst.fsm.temptari[6] ;
 wire \digitop_pav2.pie_inst.fsm.temptari[7] ;
 wire \digitop_pav2.pie_inst.fsm.temptari[8] ;
 wire \digitop_pav2.pie_inst.fsm.temptari[9] ;
 wire \digitop_pav2.pie_inst.fsm.trcal[4] ;
 wire \digitop_pav2.pie_inst.fsm.trcal[5] ;
 wire \digitop_pav2.pie_inst.fsm.trcal[6] ;
 wire \digitop_pav2.pie_inst.fsm.trcal[7] ;
 wire \digitop_pav2.pie_inst.fsm.trcal[8] ;
 wire \digitop_pav2.pie_inst.fsm.trcal[9] ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.A ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.A ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.A ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.A ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.A ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.A ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.A ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.A ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.A ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.A ;
 wire \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly10_DONT_TOUCH.A ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly10_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly11_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly12_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly13_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly14_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly15_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly16_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly17_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly18_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly19_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly1_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly20_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly21_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly22_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly23_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly24_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly2_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly3_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly4_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly5_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly6_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly7_DONT_TOUCH.Y ;
 wire \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly8_DONT_TOUCH.Y ;
 wire \digitop_pav2.proc_ctrl_inst.blf_abort ;
 wire \digitop_pav2.proc_ctrl_inst.cmd.g_sec_auth_o ;
 wire \digitop_pav2.proc_ctrl_inst.cmd.rst_b_i ;
 wire \digitop_pav2.proc_ctrl_inst.cmd.state[0] ;
 wire \digitop_pav2.proc_ctrl_inst.cmd.state[1] ;
 wire \digitop_pav2.proc_ctrl_inst.cmd.state[2] ;
 wire \digitop_pav2.proc_ctrl_inst.cmd.state[3] ;
 wire \digitop_pav2.proc_ctrl_inst.cmd.state[4] ;
 wire \digitop_pav2.proc_ctrl_inst.cmd.state[5] ;
 wire \digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[0] ;
 wire \digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[1] ;
 wire \digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[2] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.cmdctr_end3 ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.ctr[0] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.ctr[1] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.ctr[2] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.ctr[3] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.ctr[4] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.ctr[5] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.ctr[6] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.ctr[7] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.par1_en_ff ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.par2_en_ff ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.par3_en_ff ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.par4_en_ff ;
 wire \digitop_pav2.proc_ctrl_inst.cmdctr.pro_abort_b_i ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.cg_en_13 ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.cg_en_out1 ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.cg_en_out2 ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.cmd_abort_b ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_cgen.en_g_sec_i ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_cgen.fg_tc_rx_i ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate1.ck_out ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate1.w_nor ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate2.ck_out ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate2.w_nor ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.ebv_en ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.ebv_rst_b ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.fm0x_dt_tx_st_i ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.fm0x_mod_en_i ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.mode ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.n_crc_eval ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.n_pass_t1_i ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.n_rn_en ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.n_rn_rst_b ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.pass_t1_i ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.piex_dt_rx_done ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.query_dr ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.query_m[0] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.query_m[1] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.query_trext ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.rn_en ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.rn_rst_b ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[0] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[11] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[12] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[13] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[1] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[2] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[3] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[4] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[5] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[6] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[7] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[8] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.state[9] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.timeout_en_t1 ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[0] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[1] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[2] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[3] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[4] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[5] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[6] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[7] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[8] ;
 wire \digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[9] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.invalid ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[0] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[10] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[11] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[12] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[13] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[14] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[1] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[2] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[3] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[4] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[5] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[6] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[7] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[8] ;
 wire \digitop_pav2.proc_ctrl_inst.ebv.state[9] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.dif ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[0] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[10] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[11] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[12] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[13] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[14] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[15] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[1] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[2] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[3] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[4] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[5] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[6] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[7] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[8] ;
 wire \digitop_pav2.proc_ctrl_inst.inst_checker.state[9] ;
 wire \digitop_pav2.proc_ctrl_inst.int_pass_t2_flag ;
 wire \digitop_pav2.proc_ctrl_inst.int_timeout_t2 ;
 wire \digitop_pav2.proc_ctrl_inst.profsm.n_blf_abort ;
 wire \digitop_pav2.proc_ctrl_inst.profsm.r1_ff ;
 wire \digitop_pav2.proc_ctrl_inst.profsm.r1_rise_ff ;
 wire \digitop_pav2.proc_ctrl_inst.profsm.skip_abort ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_0.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_1.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_2.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_3.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_4.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_5.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_6.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_7.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_8.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_9.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_0.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_1.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_2.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_3.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_4.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_5.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_6.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_7.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_8.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_0.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_1.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_2.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_3.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_4.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_5.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_6.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_7.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_8.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_0.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_1.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_2.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_3.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_4.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_5.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_6.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_7.Y ;
 wire \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_8.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[0] ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[1] ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[2] ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[3] ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[4] ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[0] ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[1] ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[2] ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[3] ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[4] ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.pass_t2 ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.pass_t2_flag ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.ctr.piex_dt_rx_en_i ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_0.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_1.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_2.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_3.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_4.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_5.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_6.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_7.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_8.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_0.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_1.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_2.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_3.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_4.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_5.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_6.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_7.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_8.Y ;
 wire \digitop_pav2.proc_ctrl_inst.timeout.t2.jalido ;
 wire \digitop_pav2.rng_inst.rng_prngx_pav2.rngx_sec_req_i ;
 wire \digitop_pav2.rng_inst.rng_prngx_pav2.sel[0] ;
 wire \digitop_pav2.rng_inst.rng_prngx_pav2.sel[1] ;
 wire \digitop_pav2.rng_inst.rng_prngx_pav2.sel[2] ;
 wire \digitop_pav2.rng_inst.rng_prngx_pav2.trngx_data_i ;
 wire \digitop_pav2.rng_inst.rng_trngx_pav2.ff1 ;
 wire \digitop_pav2.rng_inst.rng_trngx_pav2.neg_data ;
 wire \digitop_pav2.rng_inst.rng_trngx_pav2.pos_data ;
 wire \digitop_pav2.rng_inst.rng_trngx_pav2.rngx_trngx_DONT_TOUCH.neg_data_nc ;
 wire \digitop_pav2.rng_inst.rng_trngx_pav2.xor_data ;
 wire \digitop_pav2.s1_i ;
 wire \digitop_pav2.s2_i ;
 wire \digitop_pav2.s3_i ;
 wire \digitop_pav2.sec_inst.dg_key.en_i ;
 wire \digitop_pav2.sec_inst.en_ld_data ;
 wire \digitop_pav2.sec_inst.en_ld_r ;
 wire \digitop_pav2.sec_inst.en_reg128 ;
 wire \digitop_pav2.sec_inst.en_shifto ;
 wire \digitop_pav2.sec_inst.ld_mem.round_i ;
 wire \digitop_pav2.sec_inst.ld_mem.st[0] ;
 wire \digitop_pav2.sec_inst.ld_mem.st[1] ;
 wire \digitop_pav2.sec_inst.ld_mem.st[2] ;
 wire \digitop_pav2.sec_inst.ld_mem.st[3] ;
 wire \digitop_pav2.sec_inst.ld_mem.wctr[0] ;
 wire \digitop_pav2.sec_inst.ld_mem.wctr[1] ;
 wire \digitop_pav2.sec_inst.ld_mem.wctr[2] ;
 wire \digitop_pav2.sec_inst.ld_mem.wctr[3] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[14] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[15] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[22] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[23] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[30] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[31] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[38] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[39] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[46] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[47] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[54] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[55] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[62] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[63] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[6] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[70] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[71] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[78] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[79] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[7] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[86] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[87] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[94] ;
 wire \digitop_pav2.sec_inst.ld_r.reg96_i[95] ;
 wire \digitop_pav2.sec_inst.ld_r.st[0] ;
 wire \digitop_pav2.sec_inst.ld_r.st[1] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[0] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[100] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[101] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[102] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[103] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[104] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[105] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[106] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[107] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[108] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[109] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[10] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[110] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[111] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[112] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[113] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[114] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[115] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[116] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[117] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[118] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[119] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[11] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[120] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[121] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[122] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[123] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[124] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[125] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[126] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[127] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[12] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[13] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[14] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[15] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[16] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[17] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[18] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[19] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[1] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[20] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[21] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[22] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[23] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[24] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[25] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[26] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[27] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[28] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[29] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[2] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[30] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[31] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[32] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[33] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[34] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[35] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[36] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[37] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[38] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[39] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[3] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[40] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[41] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[42] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[43] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[44] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[45] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[46] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[47] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[48] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[49] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[4] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[50] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[51] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[52] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[53] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[54] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[55] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[56] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[57] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[58] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[59] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[5] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[60] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[61] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[62] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[63] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[64] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[65] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[66] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[67] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[68] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[69] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[6] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[70] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[71] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[72] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[73] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[74] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[75] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[76] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[77] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[78] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[79] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[7] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[80] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[81] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[82] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[83] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[84] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[85] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[86] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[87] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[88] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[89] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[8] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[90] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[91] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[92] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[93] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[94] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[95] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[96] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[97] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[98] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[99] ;
 wire \digitop_pav2.sec_inst.r128.reg128_o[9] ;
 wire \digitop_pav2.sec_inst.reg160[0] ;
 wire \digitop_pav2.sec_inst.reg160[10] ;
 wire \digitop_pav2.sec_inst.reg160[11] ;
 wire \digitop_pav2.sec_inst.reg160[12] ;
 wire \digitop_pav2.sec_inst.reg160[13] ;
 wire \digitop_pav2.sec_inst.reg160[14] ;
 wire \digitop_pav2.sec_inst.reg160[15] ;
 wire \digitop_pav2.sec_inst.reg160[16] ;
 wire \digitop_pav2.sec_inst.reg160[17] ;
 wire \digitop_pav2.sec_inst.reg160[18] ;
 wire \digitop_pav2.sec_inst.reg160[19] ;
 wire \digitop_pav2.sec_inst.reg160[1] ;
 wire \digitop_pav2.sec_inst.reg160[20] ;
 wire \digitop_pav2.sec_inst.reg160[21] ;
 wire \digitop_pav2.sec_inst.reg160[22] ;
 wire \digitop_pav2.sec_inst.reg160[23] ;
 wire \digitop_pav2.sec_inst.reg160[24] ;
 wire \digitop_pav2.sec_inst.reg160[25] ;
 wire \digitop_pav2.sec_inst.reg160[26] ;
 wire \digitop_pav2.sec_inst.reg160[27] ;
 wire \digitop_pav2.sec_inst.reg160[28] ;
 wire \digitop_pav2.sec_inst.reg160[29] ;
 wire \digitop_pav2.sec_inst.reg160[2] ;
 wire \digitop_pav2.sec_inst.reg160[30] ;
 wire \digitop_pav2.sec_inst.reg160[31] ;
 wire \digitop_pav2.sec_inst.reg160[32] ;
 wire \digitop_pav2.sec_inst.reg160[33] ;
 wire \digitop_pav2.sec_inst.reg160[34] ;
 wire \digitop_pav2.sec_inst.reg160[35] ;
 wire \digitop_pav2.sec_inst.reg160[36] ;
 wire \digitop_pav2.sec_inst.reg160[37] ;
 wire \digitop_pav2.sec_inst.reg160[38] ;
 wire \digitop_pav2.sec_inst.reg160[39] ;
 wire \digitop_pav2.sec_inst.reg160[3] ;
 wire \digitop_pav2.sec_inst.reg160[40] ;
 wire \digitop_pav2.sec_inst.reg160[41] ;
 wire \digitop_pav2.sec_inst.reg160[42] ;
 wire \digitop_pav2.sec_inst.reg160[43] ;
 wire \digitop_pav2.sec_inst.reg160[44] ;
 wire \digitop_pav2.sec_inst.reg160[45] ;
 wire \digitop_pav2.sec_inst.reg160[46] ;
 wire \digitop_pav2.sec_inst.reg160[47] ;
 wire \digitop_pav2.sec_inst.reg160[48] ;
 wire \digitop_pav2.sec_inst.reg160[49] ;
 wire \digitop_pav2.sec_inst.reg160[4] ;
 wire \digitop_pav2.sec_inst.reg160[50] ;
 wire \digitop_pav2.sec_inst.reg160[51] ;
 wire \digitop_pav2.sec_inst.reg160[52] ;
 wire \digitop_pav2.sec_inst.reg160[53] ;
 wire \digitop_pav2.sec_inst.reg160[54] ;
 wire \digitop_pav2.sec_inst.reg160[55] ;
 wire \digitop_pav2.sec_inst.reg160[56] ;
 wire \digitop_pav2.sec_inst.reg160[57] ;
 wire \digitop_pav2.sec_inst.reg160[58] ;
 wire \digitop_pav2.sec_inst.reg160[59] ;
 wire \digitop_pav2.sec_inst.reg160[5] ;
 wire \digitop_pav2.sec_inst.reg160[60] ;
 wire \digitop_pav2.sec_inst.reg160[61] ;
 wire \digitop_pav2.sec_inst.reg160[62] ;
 wire \digitop_pav2.sec_inst.reg160[63] ;
 wire \digitop_pav2.sec_inst.reg160[6] ;
 wire \digitop_pav2.sec_inst.reg160[7] ;
 wire \digitop_pav2.sec_inst.reg160[8] ;
 wire \digitop_pav2.sec_inst.reg160[9] ;
 wire \digitop_pav2.sec_inst.shift_in.s1.q[0] ;
 wire \digitop_pav2.sec_inst.shift_in.s1.q[1] ;
 wire \digitop_pav2.sec_inst.shift_in.s1.q[2] ;
 wire \digitop_pav2.sec_inst.shift_in.s1.q[3] ;
 wire \digitop_pav2.sec_inst.shift_in.s1.q[4] ;
 wire \digitop_pav2.sec_inst.shift_in.s1.q[5] ;
 wire \digitop_pav2.sec_inst.shift_in.s10.q[0] ;
 wire \digitop_pav2.sec_inst.shift_in.s10.q[1] ;
 wire \digitop_pav2.sec_inst.shift_in.s10.q[2] ;
 wire \digitop_pav2.sec_inst.shift_in.s10.q[3] ;
 wire \digitop_pav2.sec_inst.shift_in.s10.q[4] ;
 wire \digitop_pav2.sec_inst.shift_in.s10.q[5] ;
 wire \digitop_pav2.sec_inst.shift_in.s11.q[0] ;
 wire \digitop_pav2.sec_inst.shift_in.s11.q[1] ;
 wire \digitop_pav2.sec_inst.shift_in.s11.q[2] ;
 wire \digitop_pav2.sec_inst.shift_in.s11.q[3] ;
 wire \digitop_pav2.sec_inst.shift_in.s11.q[4] ;
 wire \digitop_pav2.sec_inst.shift_in.s11.q[5] ;
 wire \digitop_pav2.sec_inst.shift_in.s12.q[0] ;
 wire \digitop_pav2.sec_inst.shift_in.s12.q[1] ;
 wire \digitop_pav2.sec_inst.shift_in.s12.q[2] ;
 wire \digitop_pav2.sec_inst.shift_in.s12.q[3] ;
 wire \digitop_pav2.sec_inst.shift_in.s12.q[4] ;
 wire \digitop_pav2.sec_inst.shift_in.s12.q[5] ;
 wire \digitop_pav2.sec_inst.shift_in.s2.q[0] ;
 wire \digitop_pav2.sec_inst.shift_in.s2.q[1] ;
 wire \digitop_pav2.sec_inst.shift_in.s2.q[2] ;
 wire \digitop_pav2.sec_inst.shift_in.s2.q[3] ;
 wire \digitop_pav2.sec_inst.shift_in.s2.q[4] ;
 wire \digitop_pav2.sec_inst.shift_in.s2.q[5] ;
 wire \digitop_pav2.sec_inst.shift_in.s3.q[0] ;
 wire \digitop_pav2.sec_inst.shift_in.s3.q[1] ;
 wire \digitop_pav2.sec_inst.shift_in.s3.q[2] ;
 wire \digitop_pav2.sec_inst.shift_in.s3.q[3] ;
 wire \digitop_pav2.sec_inst.shift_in.s3.q[4] ;
 wire \digitop_pav2.sec_inst.shift_in.s3.q[5] ;
 wire \digitop_pav2.sec_inst.shift_in.s4.q[0] ;
 wire \digitop_pav2.sec_inst.shift_in.s4.q[1] ;
 wire \digitop_pav2.sec_inst.shift_in.s4.q[2] ;
 wire \digitop_pav2.sec_inst.shift_in.s4.q[3] ;
 wire \digitop_pav2.sec_inst.shift_in.s4.q[4] ;
 wire \digitop_pav2.sec_inst.shift_in.s4.q[5] ;
 wire \digitop_pav2.sec_inst.shift_in.s5.q[0] ;
 wire \digitop_pav2.sec_inst.shift_in.s5.q[1] ;
 wire \digitop_pav2.sec_inst.shift_in.s5.q[2] ;
 wire \digitop_pav2.sec_inst.shift_in.s5.q[3] ;
 wire \digitop_pav2.sec_inst.shift_in.s5.q[4] ;
 wire \digitop_pav2.sec_inst.shift_in.s5.q[5] ;
 wire \digitop_pav2.sec_inst.shift_in.s6.q[0] ;
 wire \digitop_pav2.sec_inst.shift_in.s6.q[1] ;
 wire \digitop_pav2.sec_inst.shift_in.s6.q[2] ;
 wire \digitop_pav2.sec_inst.shift_in.s6.q[3] ;
 wire \digitop_pav2.sec_inst.shift_in.s6.q[4] ;
 wire \digitop_pav2.sec_inst.shift_in.s6.q[5] ;
 wire \digitop_pav2.sec_inst.shift_in.s7.q[0] ;
 wire \digitop_pav2.sec_inst.shift_in.s7.q[1] ;
 wire \digitop_pav2.sec_inst.shift_in.s7.q[2] ;
 wire \digitop_pav2.sec_inst.shift_in.s7.q[3] ;
 wire \digitop_pav2.sec_inst.shift_in.s7.q[4] ;
 wire \digitop_pav2.sec_inst.shift_in.s7.q[5] ;
 wire \digitop_pav2.sec_inst.shift_in.s8.q[0] ;
 wire \digitop_pav2.sec_inst.shift_in.s8.q[1] ;
 wire \digitop_pav2.sec_inst.shift_in.s8.q[2] ;
 wire \digitop_pav2.sec_inst.shift_in.s8.q[3] ;
 wire \digitop_pav2.sec_inst.shift_in.s8.q[4] ;
 wire \digitop_pav2.sec_inst.shift_in.s8.q[5] ;
 wire \digitop_pav2.sec_inst.shift_in.s9.q[0] ;
 wire \digitop_pav2.sec_inst.shift_in.s9.q[1] ;
 wire \digitop_pav2.sec_inst.shift_in.s9.q[2] ;
 wire \digitop_pav2.sec_inst.shift_in.s9.q[3] ;
 wire \digitop_pav2.sec_inst.shift_in.s9.q[4] ;
 wire \digitop_pav2.sec_inst.shift_in.s9.q[5] ;
 wire \digitop_pav2.sec_inst.shift_in.st[0] ;
 wire \digitop_pav2.sec_inst.shift_in.st[1] ;
 wire \digitop_pav2.sec_inst.shift_in.st[2] ;
 wire \digitop_pav2.sec_inst.shift_in.st[3] ;
 wire \digitop_pav2.sec_inst.shift_in.st[4] ;
 wire \digitop_pav2.sec_inst.shift_out.ctr[0] ;
 wire \digitop_pav2.sec_inst.shift_out.ctr[1] ;
 wire \digitop_pav2.sec_inst.shift_out.ctr[2] ;
 wire \digitop_pav2.sec_inst.shift_out.ctr[3] ;
 wire \digitop_pav2.sec_inst.shift_out.j_ctr[0] ;
 wire \digitop_pav2.sec_inst.shift_out.j_ctr[1] ;
 wire \digitop_pav2.sec_inst.shift_out.j_ctr[2] ;
 wire \digitop_pav2.sec_inst.shift_out.j_ctr[3] ;
 wire \digitop_pav2.sec_inst.shift_out.j_ctr[4] ;
 wire \digitop_pav2.sec_inst.shift_out.j_ctr[5] ;
 wire \digitop_pav2.sec_inst.shift_out.j_ctr[6] ;
 wire \digitop_pav2.sec_inst.shift_out.st[0] ;
 wire \digitop_pav2.sec_inst.shift_out.st[1] ;
 wire \digitop_pav2.sec_inst.shift_out.st[2] ;
 wire \digitop_pav2.sec_inst.shift_out.st[3] ;
 wire \digitop_pav2.sec_inst.shift_out.st[4] ;
 wire \digitop_pav2.sec_inst.shift_out.st[5] ;
 wire \digitop_pav2.sec_inst.shift_out.st[6] ;
 wire \digitop_pav2.sec_inst.shift_out.st[7] ;
 wire \digitop_pav2.sec_inst.sm.next_st[1] ;
 wire \digitop_pav2.sec_inst.sm.st[1] ;
 wire \digitop_pav2.sec_inst.sm.st[6] ;
 wire \digitop_pav2.sec_inst.sm.st[9] ;
 wire \digitop_pav2.sl_i ;
 wire \digitop_pav2.stadly_memctrl_rd_en_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt0_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt0_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt0_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt10_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt10_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt10_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt11_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt11_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt11_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt12_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt12_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt12_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt13_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt13_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt13_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt14_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt14_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt14_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt15_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt15_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt15_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt1_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt1_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt1_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt2_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt2_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt2_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt3_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt3_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt3_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt4_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt4_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt4_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt5_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt5_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt5_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt6_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt6_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt6_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt7_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt7_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt7_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt8_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt8_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt8_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt9_0.A ;
 wire \digitop_pav2.stadly_memctrl_wr_dt9_0.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_dt9_1.Y ;
 wire \digitop_pav2.stadly_memctrl_wr_en_0.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.access_clk_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.ack_clk_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.blf_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.blf_clk_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.blf_clk_pre ;
 wire \digitop_pav2.sync_inst.inst_clkx.boot_clk_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.cipher_clk_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.dft_div4_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.en_blf_fc_b ;
 wire \digitop_pav2.sync_inst.inst_clkx.fm0x_clk_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.g_access ;
 wire \digitop_pav2.sync_inst.inst_clkx.g_invent ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_fc_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_fc_clk_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_pre_clk_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_mask ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_mask_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.en_ctr ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.A ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.A ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.A ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.A ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[5].sync_pav2_clkx_delay_DONT_TOUCH.A ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[5].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.A ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[7].sync_pav2_clkx_delay_DONT_TOUCH.A ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[7].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[5].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_0.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_1.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_2.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_3.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_4.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_5.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_6.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_7.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_8.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_9.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.dis_blf_fc_b ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.en_blf_fc_b ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.mode_after_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.pass_t2_ff ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gate.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gate.w_not ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_fc_clk_gated ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_fc_clk_gated_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_gen_cg.enable ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_gen_cg.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_block_access.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_block_ack.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_block_invent.ck_out ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_block_invent.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_block_sec.ck_out ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_block_sec.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_boot.boot_dis_fix ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_boot.inst_gate.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_boot.inst_gate.w_not ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cgate.ck_in ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cgate.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cgate.w_not ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cipher.cipher_en ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cipher.inst_en.cipher_off_ff ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cipher.inst_gate.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_div_after_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_irreg_after_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_mode_after_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.cp_div_sel[0] ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.cp_div_sel[1] ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.cp_div_sel_0_after_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.cp_div_sel_1_after_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.div_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.int_rst_b ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.m2_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.m2_clk_after_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.m4_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.m4_clk_after_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.m8_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_cp.m8_clk_after_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_div4.div_gated_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_div4.div_gated_clk_before_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.div2 ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.div2_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.div4 ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div4_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div4_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_gate.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_gate.w_not ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_fm0x.en_fm0x_clk_b ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_fm0x.inst_gate.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_fm0x.inst_gate.w_not ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_ff ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_ff2 ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_ff3 ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_i ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_mem.en_mem_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_en.merge_clk_i ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_gate.ck_out ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_gate.w_or ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_merge.merge_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_piex.clkx_piex_clk_o ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_en.piex_clk_dis ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_en.slow_clk_en_b_ff2_i ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_en.slow_clk_en_b_ff3 ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_ff.slow_clk_en_b_ff ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_ff.slow_clk_en_b_i ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.enable ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.w_not ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.boot_dis_clk_after_buf ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.en_pup_clk_b ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.en_scwend_clk_b ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.en_pup_clk_b_aux ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[0] ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[1] ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[2] ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[3] ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[4] ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[5] ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.rngx_pup_clk_i ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.scwend_clk_i ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.slow_clk_en ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.trigger_clk_i ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.ck_out ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.w_not ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.ck_out ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.w_not ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_gate.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_gate.w_not ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_sel.rngx_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_trigger.trigger_clk ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.ck_out ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.w_nor ;
 wire \digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.w_not ;
 wire \digitop_pav2.sync_inst.inst_rstx.gray_counter[0] ;
 wire \digitop_pav2.sync_inst.inst_rstx.gray_counter[1] ;
 wire \digitop_pav2.sync_inst.inst_rstx.gray_counter[2] ;
 wire \digitop_pav2.sync_inst.inst_rstx.osc_clk_gated ;
 wire \digitop_pav2.sync_inst.inst_rstx.sync_rstx_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ;
 wire \digitop_pav2.sync_inst.inst_rstx.sync_rstx_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ;
 wire \digitop_pav2.sync_inst.inst_rstx.sync_rstx_gate.w_nor ;
 wire \digitop_pav2.sync_inst.inst_rstx.sync_rstx_gate.w_not ;
 wire \digitop_pav2.sync_inst.inst_rstx.trigger_DONT_TOUCH1.Q ;
 wire \digitop_pav2.testctrl_pav2.inst_enter.tm_enter ;
 wire \digitop_pav2.testctrl_pav2.inst_enter.tmrboot_clk ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[4] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[5] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[6] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[7] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[8] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[9] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.form_end ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rd_end_i ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rd_stb ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[10] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[11] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[12] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[13] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[14] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[15] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[4] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[5] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[6] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[7] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[8] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[9] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_bit ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_end_i ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_stb ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_form_enable ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_form_end ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_int_rd_stb ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_int_wr_bit ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_int_wr_stb ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.read_after_prog_ok ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[4] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[5] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[6] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[7] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[8] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[4] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[4] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[4] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[5] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_int_rd_end ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_int_wr_end ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_erase ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_prog ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_read ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_state[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.rr_erase ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.rr_prog ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.rr_read ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[4] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.int_rd_stb ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.int_wr_bit ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.int_wr_stb ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.mbist_end ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.mbist_result ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.n_int_rd_stb ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.n_int_wr_bit ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.n_int_wr_stb ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[4] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[5] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[6] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[7] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[8] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[4] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.reg_wr_en ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[4] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[5] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[6] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[7] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[8] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[9] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mbform.inst_type.tm_mbist_i ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_state[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_state[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_state[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_state[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_state[4] ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_tm_anafunc ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_tm_calclk ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_tm_clkout ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_tm_digfunc ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_tm_dummy ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_tm_mbist ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_tm_probe ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.n_tm_rnclkout ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.state[0] ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.state[1] ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.state[2] ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.state[3] ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.state[4] ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.tm_amux ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.tm_anafunc ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.tm_clkout ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.tm_digfunc ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.tm_dummy ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.tm_probe ;
 wire \digitop_pav2.testctrl_pav2.inst_mode.tm_rnclkout ;
 wire \digitop_pav2.testctrl_pav2.inst_tmamux.data_tclk_is_data ;
 wire \digitop_pav2.testctrl_pav2.inst_tmamux.window_ibias ;
 wire \digitop_pav2.testctrl_pav2.inst_tmamux.window_vcc ;
 wire \digitop_pav2.testctrl_pav2.inst_tmamux.window_vdd ;
 wire \digitop_pav2.testctrl_pav2.inst_tmamux.window_vref ;
 wire ff_erase;
 wire ff_erase_after_buf;
 wire ff_erase_ff;
 wire ff_erase_ff2;
 wire ff_erase_ff3;
 wire ff_erase_rise;
 wire ff_prog;
 wire ff_prog_after_buf;
 wire ff_prog_ff;
 wire ff_prog_ff2;
 wire ff_prog_ff3;
 wire ff_prog_rise;
 wire s1_rst_after_buf;
 wire s1_rst_ff;
 wire s1_rst_ff2;
 wire s1_set_after_buf;
 wire s1_set_ff;
 wire s1_set_ff2;
 wire s2_rst_after_buf;
 wire s2_rst_ff;
 wire s2_rst_ff2;
 wire s2_set_after_buf;
 wire s2_set_ff;
 wire s2_set_ff2;
 wire s3_rst_after_buf;
 wire s3_rst_ff;
 wire s3_rst_ff2;
 wire s3_set_after_buf;
 wire s3_set_ff;
 wire s3_set_ff2;
 wire sl_rst_after_buf;
 wire sl_rst_ff;
 wire sl_rst_ff2;
 wire sl_set_after_buf;
 wire sl_set_ff;
 wire sl_set_ff2;
 wire \stadly_mpw03_erase_rise_0.Y ;
 wire \stadly_mpw03_erase_rise_1.Y ;
 wire \stadly_mpw03_erase_rise_2.Y ;
 wire \stadly_mpw03_erase_rise_3.Y ;
 wire \stadly_mpw03_erase_rise_4.Y ;
 wire \stadly_mpw03_erase_rise_5.Y ;
 wire \stadly_mpw03_erase_rise_6.Y ;
 wire \stadly_mpw03_erase_rise_7.Y ;
 wire \stadly_mpw03_erase_rise_8.Y ;
 wire \stadly_mpw03_erase_rise_9.Y ;
 wire \stadly_mpw03_prog_rise_0.Y ;
 wire \stadly_mpw03_prog_rise_1.Y ;
 wire \stadly_mpw03_prog_rise_2.Y ;
 wire \stadly_mpw03_prog_rise_3.Y ;
 wire \stadly_mpw03_prog_rise_4.Y ;
 wire \stadly_mpw03_prog_rise_5.Y ;
 wire \stadly_mpw03_prog_rise_6.Y ;
 wire \stadly_mpw03_prog_rise_7.Y ;
 wire \stadly_mpw03_prog_rise_8.Y ;
 wire \stadly_mpw03_prog_rise_9.Y ;
 wire \vmem[0] ;
 wire \vmem[100] ;
 wire \vmem[101] ;
 wire \vmem[102] ;
 wire \vmem[103] ;
 wire \vmem[104] ;
 wire \vmem[105] ;
 wire \vmem[106] ;
 wire \vmem[107] ;
 wire \vmem[108] ;
 wire \vmem[109] ;
 wire \vmem[10] ;
 wire \vmem[110] ;
 wire \vmem[111] ;
 wire \vmem[112] ;
 wire \vmem[113] ;
 wire \vmem[114] ;
 wire \vmem[115] ;
 wire \vmem[116] ;
 wire \vmem[117] ;
 wire \vmem[118] ;
 wire \vmem[119] ;
 wire \vmem[11] ;
 wire \vmem[120] ;
 wire \vmem[121] ;
 wire \vmem[122] ;
 wire \vmem[123] ;
 wire \vmem[124] ;
 wire \vmem[125] ;
 wire \vmem[126] ;
 wire \vmem[127] ;
 wire \vmem[128] ;
 wire \vmem[129] ;
 wire \vmem[12] ;
 wire \vmem[130] ;
 wire \vmem[131] ;
 wire \vmem[132] ;
 wire \vmem[133] ;
 wire \vmem[134] ;
 wire \vmem[135] ;
 wire \vmem[136] ;
 wire \vmem[137] ;
 wire \vmem[138] ;
 wire \vmem[139] ;
 wire \vmem[13] ;
 wire \vmem[140] ;
 wire \vmem[141] ;
 wire \vmem[142] ;
 wire \vmem[143] ;
 wire \vmem[144] ;
 wire \vmem[145] ;
 wire \vmem[146] ;
 wire \vmem[147] ;
 wire \vmem[148] ;
 wire \vmem[149] ;
 wire \vmem[14] ;
 wire \vmem[150] ;
 wire \vmem[151] ;
 wire \vmem[152] ;
 wire \vmem[153] ;
 wire \vmem[154] ;
 wire \vmem[155] ;
 wire \vmem[156] ;
 wire \vmem[157] ;
 wire \vmem[158] ;
 wire \vmem[159] ;
 wire \vmem[15] ;
 wire \vmem[160] ;
 wire \vmem[161] ;
 wire \vmem[162] ;
 wire \vmem[163] ;
 wire \vmem[164] ;
 wire \vmem[165] ;
 wire \vmem[166] ;
 wire \vmem[167] ;
 wire \vmem[168] ;
 wire \vmem[169] ;
 wire \vmem[16] ;
 wire \vmem[170] ;
 wire \vmem[171] ;
 wire \vmem[172] ;
 wire \vmem[173] ;
 wire \vmem[174] ;
 wire \vmem[175] ;
 wire \vmem[176] ;
 wire \vmem[177] ;
 wire \vmem[178] ;
 wire \vmem[179] ;
 wire \vmem[17] ;
 wire \vmem[180] ;
 wire \vmem[181] ;
 wire \vmem[182] ;
 wire \vmem[183] ;
 wire \vmem[184] ;
 wire \vmem[185] ;
 wire \vmem[186] ;
 wire \vmem[187] ;
 wire \vmem[188] ;
 wire \vmem[189] ;
 wire \vmem[18] ;
 wire \vmem[190] ;
 wire \vmem[191] ;
 wire \vmem[192] ;
 wire \vmem[193] ;
 wire \vmem[194] ;
 wire \vmem[195] ;
 wire \vmem[196] ;
 wire \vmem[197] ;
 wire \vmem[198] ;
 wire \vmem[199] ;
 wire \vmem[19] ;
 wire \vmem[1] ;
 wire \vmem[200] ;
 wire \vmem[201] ;
 wire \vmem[202] ;
 wire \vmem[203] ;
 wire \vmem[204] ;
 wire \vmem[205] ;
 wire \vmem[206] ;
 wire \vmem[207] ;
 wire \vmem[208] ;
 wire \vmem[209] ;
 wire \vmem[20] ;
 wire \vmem[210] ;
 wire \vmem[211] ;
 wire \vmem[212] ;
 wire \vmem[213] ;
 wire \vmem[214] ;
 wire \vmem[215] ;
 wire \vmem[216] ;
 wire \vmem[217] ;
 wire \vmem[218] ;
 wire \vmem[219] ;
 wire \vmem[21] ;
 wire \vmem[220] ;
 wire \vmem[221] ;
 wire \vmem[222] ;
 wire \vmem[223] ;
 wire \vmem[224] ;
 wire \vmem[225] ;
 wire \vmem[226] ;
 wire \vmem[227] ;
 wire \vmem[228] ;
 wire \vmem[229] ;
 wire \vmem[22] ;
 wire \vmem[230] ;
 wire \vmem[231] ;
 wire \vmem[232] ;
 wire \vmem[233] ;
 wire \vmem[234] ;
 wire \vmem[235] ;
 wire \vmem[236] ;
 wire \vmem[237] ;
 wire \vmem[238] ;
 wire \vmem[239] ;
 wire \vmem[23] ;
 wire \vmem[240] ;
 wire \vmem[241] ;
 wire \vmem[242] ;
 wire \vmem[243] ;
 wire \vmem[244] ;
 wire \vmem[245] ;
 wire \vmem[246] ;
 wire \vmem[247] ;
 wire \vmem[248] ;
 wire \vmem[249] ;
 wire \vmem[24] ;
 wire \vmem[250] ;
 wire \vmem[251] ;
 wire \vmem[252] ;
 wire \vmem[253] ;
 wire \vmem[254] ;
 wire \vmem[255] ;
 wire \vmem[256] ;
 wire \vmem[257] ;
 wire \vmem[258] ;
 wire \vmem[259] ;
 wire \vmem[25] ;
 wire \vmem[260] ;
 wire \vmem[261] ;
 wire \vmem[262] ;
 wire \vmem[263] ;
 wire \vmem[264] ;
 wire \vmem[265] ;
 wire \vmem[266] ;
 wire \vmem[267] ;
 wire \vmem[268] ;
 wire \vmem[269] ;
 wire \vmem[26] ;
 wire \vmem[270] ;
 wire \vmem[271] ;
 wire \vmem[272] ;
 wire \vmem[273] ;
 wire \vmem[274] ;
 wire \vmem[275] ;
 wire \vmem[276] ;
 wire \vmem[277] ;
 wire \vmem[278] ;
 wire \vmem[279] ;
 wire \vmem[27] ;
 wire \vmem[280] ;
 wire \vmem[281] ;
 wire \vmem[282] ;
 wire \vmem[283] ;
 wire \vmem[284] ;
 wire \vmem[285] ;
 wire \vmem[286] ;
 wire \vmem[287] ;
 wire \vmem[288] ;
 wire \vmem[289] ;
 wire \vmem[28] ;
 wire \vmem[290] ;
 wire \vmem[291] ;
 wire \vmem[292] ;
 wire \vmem[293] ;
 wire \vmem[294] ;
 wire \vmem[295] ;
 wire \vmem[296] ;
 wire \vmem[297] ;
 wire \vmem[298] ;
 wire \vmem[299] ;
 wire \vmem[29] ;
 wire \vmem[2] ;
 wire \vmem[300] ;
 wire \vmem[301] ;
 wire \vmem[302] ;
 wire \vmem[303] ;
 wire \vmem[304] ;
 wire \vmem[305] ;
 wire \vmem[306] ;
 wire \vmem[307] ;
 wire \vmem[308] ;
 wire \vmem[309] ;
 wire \vmem[30] ;
 wire \vmem[310] ;
 wire \vmem[311] ;
 wire \vmem[312] ;
 wire \vmem[313] ;
 wire \vmem[314] ;
 wire \vmem[315] ;
 wire \vmem[316] ;
 wire \vmem[317] ;
 wire \vmem[318] ;
 wire \vmem[319] ;
 wire \vmem[31] ;
 wire \vmem[320] ;
 wire \vmem[321] ;
 wire \vmem[322] ;
 wire \vmem[323] ;
 wire \vmem[324] ;
 wire \vmem[325] ;
 wire \vmem[326] ;
 wire \vmem[327] ;
 wire \vmem[328] ;
 wire \vmem[329] ;
 wire \vmem[32] ;
 wire \vmem[330] ;
 wire \vmem[331] ;
 wire \vmem[332] ;
 wire \vmem[333] ;
 wire \vmem[334] ;
 wire \vmem[335] ;
 wire \vmem[336] ;
 wire \vmem[337] ;
 wire \vmem[338] ;
 wire \vmem[339] ;
 wire \vmem[33] ;
 wire \vmem[340] ;
 wire \vmem[341] ;
 wire \vmem[342] ;
 wire \vmem[343] ;
 wire \vmem[344] ;
 wire \vmem[345] ;
 wire \vmem[346] ;
 wire \vmem[347] ;
 wire \vmem[348] ;
 wire \vmem[349] ;
 wire \vmem[34] ;
 wire \vmem[350] ;
 wire \vmem[351] ;
 wire \vmem[352] ;
 wire \vmem[353] ;
 wire \vmem[354] ;
 wire \vmem[355] ;
 wire \vmem[356] ;
 wire \vmem[357] ;
 wire \vmem[358] ;
 wire \vmem[359] ;
 wire \vmem[35] ;
 wire \vmem[360] ;
 wire \vmem[361] ;
 wire \vmem[362] ;
 wire \vmem[363] ;
 wire \vmem[364] ;
 wire \vmem[365] ;
 wire \vmem[366] ;
 wire \vmem[367] ;
 wire \vmem[368] ;
 wire \vmem[369] ;
 wire \vmem[36] ;
 wire \vmem[370] ;
 wire \vmem[371] ;
 wire \vmem[372] ;
 wire \vmem[373] ;
 wire \vmem[374] ;
 wire \vmem[375] ;
 wire \vmem[376] ;
 wire \vmem[377] ;
 wire \vmem[378] ;
 wire \vmem[379] ;
 wire \vmem[37] ;
 wire \vmem[380] ;
 wire \vmem[381] ;
 wire \vmem[382] ;
 wire \vmem[383] ;
 wire \vmem[384] ;
 wire \vmem[385] ;
 wire \vmem[386] ;
 wire \vmem[387] ;
 wire \vmem[388] ;
 wire \vmem[389] ;
 wire \vmem[38] ;
 wire \vmem[390] ;
 wire \vmem[391] ;
 wire \vmem[392] ;
 wire \vmem[393] ;
 wire \vmem[394] ;
 wire \vmem[395] ;
 wire \vmem[396] ;
 wire \vmem[397] ;
 wire \vmem[398] ;
 wire \vmem[399] ;
 wire \vmem[39] ;
 wire \vmem[3] ;
 wire \vmem[400] ;
 wire \vmem[401] ;
 wire \vmem[402] ;
 wire \vmem[403] ;
 wire \vmem[404] ;
 wire \vmem[405] ;
 wire \vmem[406] ;
 wire \vmem[407] ;
 wire \vmem[408] ;
 wire \vmem[409] ;
 wire \vmem[40] ;
 wire \vmem[410] ;
 wire \vmem[411] ;
 wire \vmem[412] ;
 wire \vmem[413] ;
 wire \vmem[414] ;
 wire \vmem[415] ;
 wire \vmem[416] ;
 wire \vmem[417] ;
 wire \vmem[418] ;
 wire \vmem[419] ;
 wire \vmem[41] ;
 wire \vmem[420] ;
 wire \vmem[421] ;
 wire \vmem[422] ;
 wire \vmem[423] ;
 wire \vmem[424] ;
 wire \vmem[425] ;
 wire \vmem[426] ;
 wire \vmem[427] ;
 wire \vmem[428] ;
 wire \vmem[429] ;
 wire \vmem[42] ;
 wire \vmem[430] ;
 wire \vmem[431] ;
 wire \vmem[432] ;
 wire \vmem[433] ;
 wire \vmem[434] ;
 wire \vmem[435] ;
 wire \vmem[436] ;
 wire \vmem[437] ;
 wire \vmem[438] ;
 wire \vmem[439] ;
 wire \vmem[43] ;
 wire \vmem[440] ;
 wire \vmem[441] ;
 wire \vmem[442] ;
 wire \vmem[443] ;
 wire \vmem[444] ;
 wire \vmem[445] ;
 wire \vmem[446] ;
 wire \vmem[447] ;
 wire \vmem[448] ;
 wire \vmem[449] ;
 wire \vmem[44] ;
 wire \vmem[450] ;
 wire \vmem[451] ;
 wire \vmem[452] ;
 wire \vmem[453] ;
 wire \vmem[454] ;
 wire \vmem[455] ;
 wire \vmem[456] ;
 wire \vmem[457] ;
 wire \vmem[458] ;
 wire \vmem[459] ;
 wire \vmem[45] ;
 wire \vmem[460] ;
 wire \vmem[461] ;
 wire \vmem[462] ;
 wire \vmem[463] ;
 wire \vmem[464] ;
 wire \vmem[465] ;
 wire \vmem[466] ;
 wire \vmem[467] ;
 wire \vmem[468] ;
 wire \vmem[469] ;
 wire \vmem[46] ;
 wire \vmem[470] ;
 wire \vmem[471] ;
 wire \vmem[472] ;
 wire \vmem[473] ;
 wire \vmem[474] ;
 wire \vmem[475] ;
 wire \vmem[476] ;
 wire \vmem[477] ;
 wire \vmem[478] ;
 wire \vmem[479] ;
 wire \vmem[47] ;
 wire \vmem[480] ;
 wire \vmem[481] ;
 wire \vmem[482] ;
 wire \vmem[483] ;
 wire \vmem[484] ;
 wire \vmem[485] ;
 wire \vmem[486] ;
 wire \vmem[487] ;
 wire \vmem[488] ;
 wire \vmem[489] ;
 wire \vmem[48] ;
 wire \vmem[490] ;
 wire \vmem[491] ;
 wire \vmem[492] ;
 wire \vmem[493] ;
 wire \vmem[494] ;
 wire \vmem[495] ;
 wire \vmem[496] ;
 wire \vmem[497] ;
 wire \vmem[498] ;
 wire \vmem[499] ;
 wire \vmem[49] ;
 wire \vmem[4] ;
 wire \vmem[500] ;
 wire \vmem[501] ;
 wire \vmem[502] ;
 wire \vmem[503] ;
 wire \vmem[504] ;
 wire \vmem[505] ;
 wire \vmem[506] ;
 wire \vmem[507] ;
 wire \vmem[508] ;
 wire \vmem[509] ;
 wire \vmem[50] ;
 wire \vmem[510] ;
 wire \vmem[511] ;
 wire \vmem[51] ;
 wire \vmem[52] ;
 wire \vmem[53] ;
 wire \vmem[54] ;
 wire \vmem[55] ;
 wire \vmem[56] ;
 wire \vmem[57] ;
 wire \vmem[58] ;
 wire \vmem[59] ;
 wire \vmem[5] ;
 wire \vmem[60] ;
 wire \vmem[61] ;
 wire \vmem[62] ;
 wire \vmem[63] ;
 wire \vmem[64] ;
 wire \vmem[65] ;
 wire \vmem[66] ;
 wire \vmem[67] ;
 wire \vmem[68] ;
 wire \vmem[69] ;
 wire \vmem[6] ;
 wire \vmem[70] ;
 wire \vmem[71] ;
 wire \vmem[72] ;
 wire \vmem[73] ;
 wire \vmem[74] ;
 wire \vmem[75] ;
 wire \vmem[76] ;
 wire \vmem[77] ;
 wire \vmem[78] ;
 wire \vmem[79] ;
 wire \vmem[7] ;
 wire \vmem[80] ;
 wire \vmem[81] ;
 wire \vmem[82] ;
 wire \vmem[83] ;
 wire \vmem[84] ;
 wire \vmem[85] ;
 wire \vmem[86] ;
 wire \vmem[87] ;
 wire \vmem[88] ;
 wire \vmem[89] ;
 wire \vmem[8] ;
 wire \vmem[90] ;
 wire \vmem[91] ;
 wire \vmem[92] ;
 wire \vmem[93] ;
 wire \vmem[94] ;
 wire \vmem[95] ;
 wire \vmem[96] ;
 wire \vmem[97] ;
 wire \vmem[98] ;
 wire \vmem[99] ;
 wire \vmem[9] ;
 wire \vmem_after_buf[0] ;
 wire \vmem_after_buf[100] ;
 wire \vmem_after_buf[101] ;
 wire \vmem_after_buf[102] ;
 wire \vmem_after_buf[103] ;
 wire \vmem_after_buf[104] ;
 wire \vmem_after_buf[105] ;
 wire \vmem_after_buf[106] ;
 wire \vmem_after_buf[107] ;
 wire \vmem_after_buf[108] ;
 wire \vmem_after_buf[109] ;
 wire \vmem_after_buf[10] ;
 wire \vmem_after_buf[110] ;
 wire \vmem_after_buf[111] ;
 wire \vmem_after_buf[112] ;
 wire \vmem_after_buf[113] ;
 wire \vmem_after_buf[114] ;
 wire \vmem_after_buf[115] ;
 wire \vmem_after_buf[116] ;
 wire \vmem_after_buf[117] ;
 wire \vmem_after_buf[118] ;
 wire \vmem_after_buf[119] ;
 wire \vmem_after_buf[11] ;
 wire \vmem_after_buf[120] ;
 wire \vmem_after_buf[121] ;
 wire \vmem_after_buf[122] ;
 wire \vmem_after_buf[123] ;
 wire \vmem_after_buf[124] ;
 wire \vmem_after_buf[125] ;
 wire \vmem_after_buf[126] ;
 wire \vmem_after_buf[127] ;
 wire \vmem_after_buf[128] ;
 wire \vmem_after_buf[129] ;
 wire \vmem_after_buf[12] ;
 wire \vmem_after_buf[130] ;
 wire \vmem_after_buf[131] ;
 wire \vmem_after_buf[132] ;
 wire \vmem_after_buf[133] ;
 wire \vmem_after_buf[134] ;
 wire \vmem_after_buf[135] ;
 wire \vmem_after_buf[136] ;
 wire \vmem_after_buf[137] ;
 wire \vmem_after_buf[138] ;
 wire \vmem_after_buf[139] ;
 wire \vmem_after_buf[13] ;
 wire \vmem_after_buf[140] ;
 wire \vmem_after_buf[141] ;
 wire \vmem_after_buf[142] ;
 wire \vmem_after_buf[143] ;
 wire \vmem_after_buf[144] ;
 wire \vmem_after_buf[145] ;
 wire \vmem_after_buf[146] ;
 wire \vmem_after_buf[147] ;
 wire \vmem_after_buf[148] ;
 wire \vmem_after_buf[149] ;
 wire \vmem_after_buf[14] ;
 wire \vmem_after_buf[150] ;
 wire \vmem_after_buf[151] ;
 wire \vmem_after_buf[152] ;
 wire \vmem_after_buf[153] ;
 wire \vmem_after_buf[154] ;
 wire \vmem_after_buf[155] ;
 wire \vmem_after_buf[156] ;
 wire \vmem_after_buf[157] ;
 wire \vmem_after_buf[158] ;
 wire \vmem_after_buf[159] ;
 wire \vmem_after_buf[15] ;
 wire \vmem_after_buf[160] ;
 wire \vmem_after_buf[161] ;
 wire \vmem_after_buf[162] ;
 wire \vmem_after_buf[163] ;
 wire \vmem_after_buf[164] ;
 wire \vmem_after_buf[165] ;
 wire \vmem_after_buf[166] ;
 wire \vmem_after_buf[167] ;
 wire \vmem_after_buf[168] ;
 wire \vmem_after_buf[169] ;
 wire \vmem_after_buf[16] ;
 wire \vmem_after_buf[170] ;
 wire \vmem_after_buf[171] ;
 wire \vmem_after_buf[172] ;
 wire \vmem_after_buf[173] ;
 wire \vmem_after_buf[174] ;
 wire \vmem_after_buf[175] ;
 wire \vmem_after_buf[176] ;
 wire \vmem_after_buf[177] ;
 wire \vmem_after_buf[178] ;
 wire \vmem_after_buf[179] ;
 wire \vmem_after_buf[17] ;
 wire \vmem_after_buf[180] ;
 wire \vmem_after_buf[181] ;
 wire \vmem_after_buf[182] ;
 wire \vmem_after_buf[183] ;
 wire \vmem_after_buf[184] ;
 wire \vmem_after_buf[185] ;
 wire \vmem_after_buf[186] ;
 wire \vmem_after_buf[187] ;
 wire \vmem_after_buf[188] ;
 wire \vmem_after_buf[189] ;
 wire \vmem_after_buf[18] ;
 wire \vmem_after_buf[190] ;
 wire \vmem_after_buf[191] ;
 wire \vmem_after_buf[192] ;
 wire \vmem_after_buf[193] ;
 wire \vmem_after_buf[194] ;
 wire \vmem_after_buf[195] ;
 wire \vmem_after_buf[196] ;
 wire \vmem_after_buf[197] ;
 wire \vmem_after_buf[198] ;
 wire \vmem_after_buf[199] ;
 wire \vmem_after_buf[19] ;
 wire \vmem_after_buf[1] ;
 wire \vmem_after_buf[200] ;
 wire \vmem_after_buf[201] ;
 wire \vmem_after_buf[202] ;
 wire \vmem_after_buf[203] ;
 wire \vmem_after_buf[204] ;
 wire \vmem_after_buf[205] ;
 wire \vmem_after_buf[206] ;
 wire \vmem_after_buf[207] ;
 wire \vmem_after_buf[208] ;
 wire \vmem_after_buf[209] ;
 wire \vmem_after_buf[20] ;
 wire \vmem_after_buf[210] ;
 wire \vmem_after_buf[211] ;
 wire \vmem_after_buf[212] ;
 wire \vmem_after_buf[213] ;
 wire \vmem_after_buf[214] ;
 wire \vmem_after_buf[215] ;
 wire \vmem_after_buf[216] ;
 wire \vmem_after_buf[217] ;
 wire \vmem_after_buf[218] ;
 wire \vmem_after_buf[219] ;
 wire \vmem_after_buf[21] ;
 wire \vmem_after_buf[220] ;
 wire \vmem_after_buf[221] ;
 wire \vmem_after_buf[222] ;
 wire \vmem_after_buf[223] ;
 wire \vmem_after_buf[224] ;
 wire \vmem_after_buf[225] ;
 wire \vmem_after_buf[226] ;
 wire \vmem_after_buf[227] ;
 wire \vmem_after_buf[228] ;
 wire \vmem_after_buf[229] ;
 wire \vmem_after_buf[22] ;
 wire \vmem_after_buf[230] ;
 wire \vmem_after_buf[231] ;
 wire \vmem_after_buf[232] ;
 wire \vmem_after_buf[233] ;
 wire \vmem_after_buf[234] ;
 wire \vmem_after_buf[235] ;
 wire \vmem_after_buf[236] ;
 wire \vmem_after_buf[237] ;
 wire \vmem_after_buf[238] ;
 wire \vmem_after_buf[239] ;
 wire \vmem_after_buf[23] ;
 wire \vmem_after_buf[240] ;
 wire \vmem_after_buf[241] ;
 wire \vmem_after_buf[242] ;
 wire \vmem_after_buf[243] ;
 wire \vmem_after_buf[244] ;
 wire \vmem_after_buf[245] ;
 wire \vmem_after_buf[246] ;
 wire \vmem_after_buf[247] ;
 wire \vmem_after_buf[248] ;
 wire \vmem_after_buf[249] ;
 wire \vmem_after_buf[24] ;
 wire \vmem_after_buf[250] ;
 wire \vmem_after_buf[251] ;
 wire \vmem_after_buf[252] ;
 wire \vmem_after_buf[253] ;
 wire \vmem_after_buf[254] ;
 wire \vmem_after_buf[255] ;
 wire \vmem_after_buf[256] ;
 wire \vmem_after_buf[257] ;
 wire \vmem_after_buf[258] ;
 wire \vmem_after_buf[259] ;
 wire \vmem_after_buf[25] ;
 wire \vmem_after_buf[260] ;
 wire \vmem_after_buf[261] ;
 wire \vmem_after_buf[262] ;
 wire \vmem_after_buf[263] ;
 wire \vmem_after_buf[264] ;
 wire \vmem_after_buf[265] ;
 wire \vmem_after_buf[266] ;
 wire \vmem_after_buf[267] ;
 wire \vmem_after_buf[268] ;
 wire \vmem_after_buf[269] ;
 wire \vmem_after_buf[26] ;
 wire \vmem_after_buf[270] ;
 wire \vmem_after_buf[271] ;
 wire \vmem_after_buf[272] ;
 wire \vmem_after_buf[273] ;
 wire \vmem_after_buf[274] ;
 wire \vmem_after_buf[275] ;
 wire \vmem_after_buf[276] ;
 wire \vmem_after_buf[277] ;
 wire \vmem_after_buf[278] ;
 wire \vmem_after_buf[279] ;
 wire \vmem_after_buf[27] ;
 wire \vmem_after_buf[280] ;
 wire \vmem_after_buf[281] ;
 wire \vmem_after_buf[282] ;
 wire \vmem_after_buf[283] ;
 wire \vmem_after_buf[284] ;
 wire \vmem_after_buf[285] ;
 wire \vmem_after_buf[286] ;
 wire \vmem_after_buf[287] ;
 wire \vmem_after_buf[288] ;
 wire \vmem_after_buf[289] ;
 wire \vmem_after_buf[28] ;
 wire \vmem_after_buf[290] ;
 wire \vmem_after_buf[291] ;
 wire \vmem_after_buf[292] ;
 wire \vmem_after_buf[293] ;
 wire \vmem_after_buf[294] ;
 wire \vmem_after_buf[295] ;
 wire \vmem_after_buf[296] ;
 wire \vmem_after_buf[297] ;
 wire \vmem_after_buf[298] ;
 wire \vmem_after_buf[299] ;
 wire \vmem_after_buf[29] ;
 wire \vmem_after_buf[2] ;
 wire \vmem_after_buf[300] ;
 wire \vmem_after_buf[301] ;
 wire \vmem_after_buf[302] ;
 wire \vmem_after_buf[303] ;
 wire \vmem_after_buf[304] ;
 wire \vmem_after_buf[305] ;
 wire \vmem_after_buf[306] ;
 wire \vmem_after_buf[307] ;
 wire \vmem_after_buf[308] ;
 wire \vmem_after_buf[309] ;
 wire \vmem_after_buf[30] ;
 wire \vmem_after_buf[310] ;
 wire \vmem_after_buf[311] ;
 wire \vmem_after_buf[312] ;
 wire \vmem_after_buf[313] ;
 wire \vmem_after_buf[314] ;
 wire \vmem_after_buf[315] ;
 wire \vmem_after_buf[316] ;
 wire \vmem_after_buf[317] ;
 wire \vmem_after_buf[318] ;
 wire \vmem_after_buf[319] ;
 wire \vmem_after_buf[31] ;
 wire \vmem_after_buf[320] ;
 wire \vmem_after_buf[321] ;
 wire \vmem_after_buf[322] ;
 wire \vmem_after_buf[323] ;
 wire \vmem_after_buf[324] ;
 wire \vmem_after_buf[325] ;
 wire \vmem_after_buf[326] ;
 wire \vmem_after_buf[327] ;
 wire \vmem_after_buf[328] ;
 wire \vmem_after_buf[329] ;
 wire \vmem_after_buf[32] ;
 wire \vmem_after_buf[330] ;
 wire \vmem_after_buf[331] ;
 wire \vmem_after_buf[332] ;
 wire \vmem_after_buf[333] ;
 wire \vmem_after_buf[334] ;
 wire \vmem_after_buf[335] ;
 wire \vmem_after_buf[336] ;
 wire \vmem_after_buf[337] ;
 wire \vmem_after_buf[338] ;
 wire \vmem_after_buf[339] ;
 wire \vmem_after_buf[33] ;
 wire \vmem_after_buf[340] ;
 wire \vmem_after_buf[341] ;
 wire \vmem_after_buf[342] ;
 wire \vmem_after_buf[343] ;
 wire \vmem_after_buf[344] ;
 wire \vmem_after_buf[345] ;
 wire \vmem_after_buf[346] ;
 wire \vmem_after_buf[347] ;
 wire \vmem_after_buf[348] ;
 wire \vmem_after_buf[349] ;
 wire \vmem_after_buf[34] ;
 wire \vmem_after_buf[350] ;
 wire \vmem_after_buf[351] ;
 wire \vmem_after_buf[352] ;
 wire \vmem_after_buf[353] ;
 wire \vmem_after_buf[354] ;
 wire \vmem_after_buf[355] ;
 wire \vmem_after_buf[356] ;
 wire \vmem_after_buf[357] ;
 wire \vmem_after_buf[358] ;
 wire \vmem_after_buf[359] ;
 wire \vmem_after_buf[35] ;
 wire \vmem_after_buf[360] ;
 wire \vmem_after_buf[361] ;
 wire \vmem_after_buf[362] ;
 wire \vmem_after_buf[363] ;
 wire \vmem_after_buf[364] ;
 wire \vmem_after_buf[365] ;
 wire \vmem_after_buf[366] ;
 wire \vmem_after_buf[367] ;
 wire \vmem_after_buf[368] ;
 wire \vmem_after_buf[369] ;
 wire \vmem_after_buf[36] ;
 wire \vmem_after_buf[370] ;
 wire \vmem_after_buf[371] ;
 wire \vmem_after_buf[372] ;
 wire \vmem_after_buf[373] ;
 wire \vmem_after_buf[374] ;
 wire \vmem_after_buf[375] ;
 wire \vmem_after_buf[376] ;
 wire \vmem_after_buf[377] ;
 wire \vmem_after_buf[378] ;
 wire \vmem_after_buf[379] ;
 wire \vmem_after_buf[37] ;
 wire \vmem_after_buf[380] ;
 wire \vmem_after_buf[381] ;
 wire \vmem_after_buf[382] ;
 wire \vmem_after_buf[383] ;
 wire \vmem_after_buf[384] ;
 wire \vmem_after_buf[385] ;
 wire \vmem_after_buf[386] ;
 wire \vmem_after_buf[387] ;
 wire \vmem_after_buf[388] ;
 wire \vmem_after_buf[389] ;
 wire \vmem_after_buf[38] ;
 wire \vmem_after_buf[390] ;
 wire \vmem_after_buf[391] ;
 wire \vmem_after_buf[392] ;
 wire \vmem_after_buf[393] ;
 wire \vmem_after_buf[394] ;
 wire \vmem_after_buf[395] ;
 wire \vmem_after_buf[396] ;
 wire \vmem_after_buf[397] ;
 wire \vmem_after_buf[398] ;
 wire \vmem_after_buf[399] ;
 wire \vmem_after_buf[39] ;
 wire \vmem_after_buf[3] ;
 wire \vmem_after_buf[400] ;
 wire \vmem_after_buf[401] ;
 wire \vmem_after_buf[402] ;
 wire \vmem_after_buf[403] ;
 wire \vmem_after_buf[404] ;
 wire \vmem_after_buf[405] ;
 wire \vmem_after_buf[406] ;
 wire \vmem_after_buf[407] ;
 wire \vmem_after_buf[408] ;
 wire \vmem_after_buf[409] ;
 wire \vmem_after_buf[40] ;
 wire \vmem_after_buf[410] ;
 wire \vmem_after_buf[411] ;
 wire \vmem_after_buf[412] ;
 wire \vmem_after_buf[413] ;
 wire \vmem_after_buf[414] ;
 wire \vmem_after_buf[415] ;
 wire \vmem_after_buf[416] ;
 wire \vmem_after_buf[417] ;
 wire \vmem_after_buf[418] ;
 wire \vmem_after_buf[419] ;
 wire \vmem_after_buf[41] ;
 wire \vmem_after_buf[420] ;
 wire \vmem_after_buf[421] ;
 wire \vmem_after_buf[422] ;
 wire \vmem_after_buf[423] ;
 wire \vmem_after_buf[424] ;
 wire \vmem_after_buf[425] ;
 wire \vmem_after_buf[426] ;
 wire \vmem_after_buf[427] ;
 wire \vmem_after_buf[428] ;
 wire \vmem_after_buf[429] ;
 wire \vmem_after_buf[42] ;
 wire \vmem_after_buf[430] ;
 wire \vmem_after_buf[431] ;
 wire \vmem_after_buf[432] ;
 wire \vmem_after_buf[433] ;
 wire \vmem_after_buf[434] ;
 wire \vmem_after_buf[435] ;
 wire \vmem_after_buf[436] ;
 wire \vmem_after_buf[437] ;
 wire \vmem_after_buf[438] ;
 wire \vmem_after_buf[439] ;
 wire \vmem_after_buf[43] ;
 wire \vmem_after_buf[440] ;
 wire \vmem_after_buf[441] ;
 wire \vmem_after_buf[442] ;
 wire \vmem_after_buf[443] ;
 wire \vmem_after_buf[444] ;
 wire \vmem_after_buf[445] ;
 wire \vmem_after_buf[446] ;
 wire \vmem_after_buf[447] ;
 wire \vmem_after_buf[448] ;
 wire \vmem_after_buf[449] ;
 wire \vmem_after_buf[44] ;
 wire \vmem_after_buf[450] ;
 wire \vmem_after_buf[451] ;
 wire \vmem_after_buf[452] ;
 wire \vmem_after_buf[453] ;
 wire \vmem_after_buf[454] ;
 wire \vmem_after_buf[455] ;
 wire \vmem_after_buf[456] ;
 wire \vmem_after_buf[457] ;
 wire \vmem_after_buf[458] ;
 wire \vmem_after_buf[459] ;
 wire \vmem_after_buf[45] ;
 wire \vmem_after_buf[460] ;
 wire \vmem_after_buf[461] ;
 wire \vmem_after_buf[462] ;
 wire \vmem_after_buf[463] ;
 wire \vmem_after_buf[464] ;
 wire \vmem_after_buf[465] ;
 wire \vmem_after_buf[466] ;
 wire \vmem_after_buf[467] ;
 wire \vmem_after_buf[468] ;
 wire \vmem_after_buf[469] ;
 wire \vmem_after_buf[46] ;
 wire \vmem_after_buf[470] ;
 wire \vmem_after_buf[471] ;
 wire \vmem_after_buf[472] ;
 wire \vmem_after_buf[473] ;
 wire \vmem_after_buf[474] ;
 wire \vmem_after_buf[475] ;
 wire \vmem_after_buf[476] ;
 wire \vmem_after_buf[477] ;
 wire \vmem_after_buf[478] ;
 wire \vmem_after_buf[479] ;
 wire \vmem_after_buf[47] ;
 wire \vmem_after_buf[480] ;
 wire \vmem_after_buf[481] ;
 wire \vmem_after_buf[482] ;
 wire \vmem_after_buf[483] ;
 wire \vmem_after_buf[484] ;
 wire \vmem_after_buf[485] ;
 wire \vmem_after_buf[486] ;
 wire \vmem_after_buf[487] ;
 wire \vmem_after_buf[488] ;
 wire \vmem_after_buf[489] ;
 wire \vmem_after_buf[48] ;
 wire \vmem_after_buf[490] ;
 wire \vmem_after_buf[491] ;
 wire \vmem_after_buf[492] ;
 wire \vmem_after_buf[493] ;
 wire \vmem_after_buf[494] ;
 wire \vmem_after_buf[495] ;
 wire \vmem_after_buf[496] ;
 wire \vmem_after_buf[497] ;
 wire \vmem_after_buf[498] ;
 wire \vmem_after_buf[499] ;
 wire \vmem_after_buf[49] ;
 wire \vmem_after_buf[4] ;
 wire \vmem_after_buf[500] ;
 wire \vmem_after_buf[501] ;
 wire \vmem_after_buf[502] ;
 wire \vmem_after_buf[503] ;
 wire \vmem_after_buf[504] ;
 wire \vmem_after_buf[505] ;
 wire \vmem_after_buf[506] ;
 wire \vmem_after_buf[507] ;
 wire \vmem_after_buf[508] ;
 wire \vmem_after_buf[509] ;
 wire \vmem_after_buf[50] ;
 wire \vmem_after_buf[510] ;
 wire \vmem_after_buf[511] ;
 wire \vmem_after_buf[51] ;
 wire \vmem_after_buf[52] ;
 wire \vmem_after_buf[53] ;
 wire \vmem_after_buf[54] ;
 wire \vmem_after_buf[55] ;
 wire \vmem_after_buf[56] ;
 wire \vmem_after_buf[57] ;
 wire \vmem_after_buf[58] ;
 wire \vmem_after_buf[59] ;
 wire \vmem_after_buf[5] ;
 wire \vmem_after_buf[60] ;
 wire \vmem_after_buf[61] ;
 wire \vmem_after_buf[62] ;
 wire \vmem_after_buf[63] ;
 wire \vmem_after_buf[64] ;
 wire \vmem_after_buf[65] ;
 wire \vmem_after_buf[66] ;
 wire \vmem_after_buf[67] ;
 wire \vmem_after_buf[68] ;
 wire \vmem_after_buf[69] ;
 wire \vmem_after_buf[6] ;
 wire \vmem_after_buf[70] ;
 wire \vmem_after_buf[71] ;
 wire \vmem_after_buf[72] ;
 wire \vmem_after_buf[73] ;
 wire \vmem_after_buf[74] ;
 wire \vmem_after_buf[75] ;
 wire \vmem_after_buf[76] ;
 wire \vmem_after_buf[77] ;
 wire \vmem_after_buf[78] ;
 wire \vmem_after_buf[79] ;
 wire \vmem_after_buf[7] ;
 wire \vmem_after_buf[80] ;
 wire \vmem_after_buf[81] ;
 wire \vmem_after_buf[82] ;
 wire \vmem_after_buf[83] ;
 wire \vmem_after_buf[84] ;
 wire \vmem_after_buf[85] ;
 wire \vmem_after_buf[86] ;
 wire \vmem_after_buf[87] ;
 wire \vmem_after_buf[88] ;
 wire \vmem_after_buf[89] ;
 wire \vmem_after_buf[8] ;
 wire \vmem_after_buf[90] ;
 wire \vmem_after_buf[91] ;
 wire \vmem_after_buf[92] ;
 wire \vmem_after_buf[93] ;
 wire \vmem_after_buf[94] ;
 wire \vmem_after_buf[95] ;
 wire \vmem_after_buf[96] ;
 wire \vmem_after_buf[97] ;
 wire \vmem_after_buf[98] ;
 wire \vmem_after_buf[99] ;
 wire \vmem_after_buf[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1609;
 wire net1616;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 inv_2 _11536_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[3] ),
    .Y(_07020_));
 inv_2 _11537_ (.A(\digitop_pav2.access_inst.access_ctrl0.proc_rd_finish_i ),
    .Y(_07021_));
 inv_2 _11538_ (.A(\digitop_pav2.access_inst.access_ctrl0.rx_par1_i ),
    .Y(_07022_));
 inv_2 _11539_ (.A(\digitop_pav2.access_inst.access_ctrl0.ld_key_env_finish_i ),
    .Y(_07023_));
 inv_2 _11540_ (.A(net1046),
    .Y(_07024_));
 inv_2 _11541_ (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[1] ),
    .Y(_07025_));
 inv_2 _11542_ (.A(net1049),
    .Y(_07026_));
 inv_2 _11543_ (.A(net1053),
    .Y(_07027_));
 inv_2 _11544_ (.A(net1056),
    .Y(_07028_));
 inv_2 _11545_ (.A(net1058),
    .Y(_07029_));
 inv_2 _11546_ (.A(net1063),
    .Y(_07030_));
 inv_2 _11547_ (.A(\digitop_pav2.access_inst.access_ctrl0.prev_busy ),
    .Y(_07031_));
 inv_2 _11548_ (.A(net1066),
    .Y(_07032_));
 inv_2 _11549_ (.A(\digitop_pav2.access_inst.access_check0.ctrl_wcknzero_ck ),
    .Y(_07033_));
 inv_2 _11550_ (.A(\digitop_pav2.access_inst.access_check0.mem_sign_check_sync_o ),
    .Y(_07034_));
 inv_2 _11551_ (.A(net1068),
    .Y(_07035_));
 inv_2 _11552_ (.A(\digitop_pav2.access_inst.access_ctrl0.dt_acc_done ),
    .Y(_07036_));
 inv_2 _11553_ (.A(\digitop_pav2.access_inst.access_ctrl0.replay_nok ),
    .Y(_07037_));
 inv_2 _11554_ (.A(\digitop_pav2.access_inst.access_ctrl0.replay_ok ),
    .Y(_07038_));
 inv_2 _11555_ (.A(net1071),
    .Y(_07039_));
 inv_2 _11556_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[1] ),
    .Y(_07040_));
 inv_2 _11557_ (.A(net1302),
    .Y(_07041_));
 inv_2 _11558_ (.A(\digitop_pav2.crc_inst.crc5_q[2] ),
    .Y(_07042_));
 inv_2 _11559_ (.A(\digitop_pav2.crc_inst.crc16_q[15] ),
    .Y(_07043_));
 inv_2 _11560_ (.A(\digitop_pav2.crc_inst.crc16_q[11] ),
    .Y(_07044_));
 inv_2 _11561_ (.A(\digitop_pav2.crc_inst.crc16_q[4] ),
    .Y(_07045_));
 inv_2 _11562_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_s_ff_i ),
    .Y(_07046_));
 inv_2 _11563_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_s_ff_i ),
    .Y(_07047_));
 inv_2 _11564_ (.A(net1251),
    .Y(_07048_));
 inv_2 _11565_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_mem.en_mem_clk ),
    .Y(_07049_));
 inv_2 _11566_ (.A(net1153),
    .Y(_07050_));
 inv_2 _11567_ (.A(net1156),
    .Y(_07051_));
 inv_2 _11568_ (.A(net1159),
    .Y(_07052_));
 inv_2 _11569_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[0] ),
    .Y(_07053_));
 inv_2 _11570_ (.A(\digitop_pav2.ack_inst.cnt_ff[0] ),
    .Y(_07054_));
 inv_2 _11571_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[0] ),
    .Y(_07055_));
 inv_2 _11572_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[0] ),
    .Y(_07056_));
 inv_2 _11573_ (.A(net1707),
    .Y(_07057_));
 inv_2 _11574_ (.A(\digitop_pav2.boot_inst.boot_ctrl0.proc_crc_end_i ),
    .Y(_07058_));
 inv_2 _11575_ (.A(\digitop_pav2.boot_inst.boot_ctrl0.proc_boot_end_i ),
    .Y(_07059_));
 inv_2 _11576_ (.A(net1446),
    .Y(_07060_));
 inv_2 _11577_ (.A(net1084),
    .Y(_07061_));
 inv_2 _11578_ (.A(\digitop_pav2.ack_inst.rcnt_ff[1] ),
    .Y(_07062_));
 inv_2 _11579_ (.A(net1691),
    .Y(_07063_));
 inv_2 _11580_ (.A(net702),
    .Y(_07064_));
 inv_2 _11581_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[5] ),
    .Y(_07065_));
 inv_2 _11582_ (.A(net1253),
    .Y(_07066_));
 inv_2 _11583_ (.A(net1254),
    .Y(_07067_));
 inv_2 _11584_ (.A(net1260),
    .Y(_07068_));
 inv_2 _11585_ (.A(net1694),
    .Y(_07069_));
 inv_2 _11586_ (.A(net1295),
    .Y(_07070_));
 inv_2 _11587_ (.A(\digitop_pav2.crc_inst.dt_rx_i ),
    .Y(_07071_));
 inv_2 _11588_ (.A(\digitop_pav2.memctrl_inst.state[0] ),
    .Y(_07072_));
 inv_2 _11589_ (.A(net1135),
    .Y(_07073_));
 inv_2 _11590_ (.A(\digitop_pav2.memctrl_inst.flops_0x081[2] ),
    .Y(_07074_));
 inv_2 _11591_ (.A(net1127),
    .Y(_07075_));
 inv_2 _11592_ (.A(net1121),
    .Y(_07076_));
 inv_2 _11593_ (.A(net1118),
    .Y(_07077_));
 inv_2 _11594_ (.A(net1117),
    .Y(_07078_));
 inv_2 _11595_ (.A(net1110),
    .Y(_07079_));
 inv_2 _11596_ (.A(net1099),
    .Y(_07080_));
 inv_2 _11597_ (.A(net1095),
    .Y(_07081_));
 inv_2 _11598_ (.A(net1093),
    .Y(_07082_));
 inv_2 _11599_ (.A(net1087),
    .Y(_07083_));
 inv_2 _11600_ (.A(net1484),
    .Y(_07084_));
 inv_2 _11601_ (.A(net1486),
    .Y(_07085_));
 inv_2 _11602_ (.A(net1650),
    .Y(_07086_));
 inv_2 _11603_ (.A(net1286),
    .Y(_07087_));
 inv_2 _11604_ (.A(\digitop_pav2.ack_inst.cnt_ff[2] ),
    .Y(_07088_));
 inv_2 _11605_ (.A(\digitop_pav2.ack_inst.cnt_ff[3] ),
    .Y(_07089_));
 inv_2 _11606_ (.A(net1142),
    .Y(_07090_));
 inv_2 _11607_ (.A(net1151),
    .Y(_07091_));
 inv_2 _11608_ (.A(net472),
    .Y(_07092_));
 inv_2 _11609_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[2] ),
    .Y(_07093_));
 inv_2 _11610_ (.A(net443),
    .Y(_07094_));
 inv_2 _11611_ (.A(\digitop_pav2.access_inst.access_check0.fg_i[1] ),
    .Y(_07095_));
 inv_2 _11612_ (.A(\digitop_pav2.access_inst.access_check0.fg_i[3] ),
    .Y(_07096_));
 inv_2 _11613_ (.A(\digitop_pav2.access_inst.access_check0.fg_i[5] ),
    .Y(_07097_));
 inv_2 _11614_ (.A(\digitop_pav2.access_inst.access_check0.fg_i[6] ),
    .Y(_07098_));
 inv_2 _11615_ (.A(\digitop_pav2.access_inst.access_check0.fg_i[7] ),
    .Y(_07099_));
 inv_2 _11616_ (.A(\digitop_pav2.boot_inst.boot_proc0.proc_mask[3] ),
    .Y(_07100_));
 inv_2 _11617_ (.A(\digitop_pav2.boot_inst.boot_proc0.proc_fg[12] ),
    .Y(_07101_));
 inv_2 _11618_ (.A(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[9] ),
    .Y(_07102_));
 inv_2 _11619_ (.A(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[13] ),
    .Y(_07103_));
 inv_2 _11620_ (.A(\digitop_pav2.access_inst.access_check0.pc_lock_check_i ),
    .Y(_07104_));
 inv_2 _11621_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[1] ),
    .Y(_07105_));
 clkinv_4 _11622_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[2] ),
    .Y(_07106_));
 inv_2 _11623_ (.A(\digitop_pav2.rng_inst.rng_prngx_pav2.rngx_sec_req_i ),
    .Y(_07107_));
 inv_2 _11624_ (.A(\digitop_pav2.sec_inst.dg_key.en_i ),
    .Y(_07108_));
 inv_2 _11625_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_9.Y ),
    .Y(_07109_));
 inv_2 _11626_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_9.Y ),
    .Y(_07110_));
 inv_2 _11627_ (.A(net970),
    .Y(_07111_));
 inv_2 _11628_ (.A(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_2b_o ),
    .Y(_07112_));
 inv_2 _11629_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.tm_digfunc ),
    .Y(_07113_));
 inv_2 _11630_ (.A(net413),
    .Y(_07114_));
 inv_2 _11631_ (.A(net1826),
    .Y(_07115_));
 inv_2 _11632_ (.A(\digitop_pav2.cal_inst.calx_mux.dtest_trim_1_i ),
    .Y(_07116_));
 inv_2 _11633_ (.A(\digitop_pav2.cal_inst.calx_mux.dtest_trim_0_i ),
    .Y(_07117_));
 inv_2 _11634_ (.A(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[3] ),
    .Y(_07118_));
 inv_2 _11635_ (.A(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[4] ),
    .Y(_07119_));
 inv_2 _11636_ (.A(net709),
    .Y(_07120_));
 inv_2 _11637_ (.A(\digitop_pav2.sec_inst.shift_out.st[0] ),
    .Y(_07121_));
 inv_2 _11638_ (.A(net188),
    .Y(_07122_));
 inv_2 _11639_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[0] ),
    .Y(_07123_));
 inv_2 _11640_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[3] ),
    .Y(_07124_));
 inv_2 _11641_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[2] ),
    .Y(_07125_));
 inv_2 _11642_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[1] ),
    .Y(_07126_));
 inv_2 _11643_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.flags_en_o ),
    .Y(_07127_));
 inv_2 _11644_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.mask_mismatch_ff ),
    .Y(_07128_));
 inv_2 _11645_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[5] ),
    .Y(_07129_));
 inv_2 _11646_ (.A(\digitop_pav2.proc_ctrl_inst.int_timeout_t2 ),
    .Y(_07130_));
 inv_2 _11647_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.select_valid_o ),
    .Y(_07131_));
 inv_2 _11648_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[7] ),
    .Y(_07132_));
 inv_2 _11649_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[6] ),
    .Y(_07133_));
 inv_2 _11650_ (.A(net1176),
    .Y(_07134_));
 inv_2 _11651_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[4] ),
    .Y(_07135_));
 inv_2 _11652_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[0] ),
    .Y(_07136_));
 inv_2 _11653_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[0] ),
    .Y(_07137_));
 inv_2 _11654_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[7] ),
    .Y(_07138_));
 inv_2 _11655_ (.A(\digitop_pav2.func_rr_read ),
    .Y(_07139_));
 inv_2 _11656_ (.A(\digitop_pav2.memctrl_inst.state[1] ),
    .Y(_07140_));
 inv_2 _11657_ (.A(\digitop_pav2.memctrl_inst.reg_wr_ok_ff2 ),
    .Y(_07141_));
 inv_2 _11658_ (.A(\digitop_pav2.stadly_memctrl_wr_dt1_1.Y ),
    .Y(_07142_));
 inv_2 _11659_ (.A(\digitop_pav2.stadly_memctrl_wr_dt2_1.Y ),
    .Y(_07143_));
 inv_2 _11660_ (.A(\digitop_pav2.stadly_memctrl_wr_dt6_1.Y ),
    .Y(_07144_));
 inv_2 _11661_ (.A(\digitop_pav2.pie_inst.fsm.state[0] ),
    .Y(_07145_));
 inv_2 _11662_ (.A(\digitop_pav2.pie_inst.fsm.dif_pos_fix[0] ),
    .Y(_07146_));
 inv_2 _11663_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[1] ),
    .Y(_07147_));
 inv_2 _11664_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[3] ),
    .Y(_07148_));
 inv_2 _11665_ (.A(\digitop_pav2.pie_inst.fsm.pivot[0] ),
    .Y(_07149_));
 inv_2 _11666_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.pass_t1_i ),
    .Y(_07150_));
 inv_2 _11667_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_end_i ),
    .Y(_07151_));
 inv_2 _11668_ (.A(net1480),
    .Y(_07152_));
 inv_2 _11669_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_cgen.fg_tc_rx_i ),
    .Y(_07153_));
 inv_2 _11670_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[2] ),
    .Y(_07154_));
 inv_2 _11671_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[5] ),
    .Y(_07155_));
 inv_2 _11672_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[3] ),
    .Y(_07156_));
 inv_2 _11673_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[3] ),
    .Y(_07157_));
 inv_2 _11674_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[4] ),
    .Y(_07158_));
 inv_2 _11675_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.en_ctr ),
    .Y(_00154_));
 inv_2 _11676_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Y(_00146_));
 inv_2 _11677_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Y(_00147_));
 inv_2 _11678_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Y(_00148_));
 inv_2 _11679_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Y(_00149_));
 inv_2 _11680_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Y(_00150_));
 inv_2 _11681_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[5].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Y(_00151_));
 inv_2 _11682_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Y(_00152_));
 inv_2 _11683_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[7].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Y(_00153_));
 inv_2 _11684_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.reg_wr_en ),
    .Y(_07159_));
 inv_2 _11685_ (.A(\digitop_pav2.proc_ctrl_inst.profsm.r1_ff ),
    .Y(_07160_));
 inv_2 _11686_ (.A(\digitop_pav2.proc_ctrl_inst.profsm.r1_rise_ff ),
    .Y(_07161_));
 inv_2 _11687_ (.A(net969),
    .Y(_07162_));
 inv_2 _11688_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.tm_amux ),
    .Y(_07163_));
 inv_2 _11689_ (.A(net711),
    .Y(_07164_));
 inv_2 _11690_ (.A(\digitop_pav2.func_rnclk_en ),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_ff.slow_clk_en_b_i ));
 inv_2 _11691_ (.A(\digitop_pav2.pie_inst.fsm.neg_i[1] ),
    .Y(_07165_));
 inv_2 _11692_ (.A(tclk_i),
    .Y(_00203_));
 inv_2 _11693_ (.A(net68),
    .Y(_07166_));
 inv_2 _11694_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.tm_anafunc ),
    .Y(_07167_));
 inv_2 _11695_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.tm_probe ),
    .Y(_07168_));
 inv_2 _11696_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.mbist_result ),
    .Y(_07169_));
 inv_2 _11697_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.t2.jalido ),
    .Y(_07170_));
 inv_2 _11698_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[8] ),
    .Y(_07171_));
 inv_2 _11699_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[8] ),
    .Y(_07172_));
 inv_2 _11700_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[9] ),
    .Y(_07173_));
 inv_2 _11701_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[9] ),
    .Y(_07174_));
 inv_2 _11702_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[10] ),
    .Y(_07175_));
 inv_2 _11703_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[10] ),
    .Y(_07176_));
 inv_2 _11704_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[11] ),
    .Y(_07177_));
 inv_2 _11705_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[11] ),
    .Y(_07178_));
 inv_2 _11706_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[12] ),
    .Y(_07179_));
 inv_2 _11707_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[12] ),
    .Y(_07180_));
 inv_2 _11708_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[13] ),
    .Y(_07181_));
 inv_2 _11709_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[13] ),
    .Y(_07182_));
 inv_2 _11710_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[14] ),
    .Y(_07183_));
 inv_2 _11711_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[14] ),
    .Y(_07184_));
 inv_2 _11712_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[15] ),
    .Y(_07185_));
 inv_2 _11713_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[15] ),
    .Y(_07186_));
 inv_2 _11714_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[8] ),
    .Y(_07187_));
 inv_2 _11715_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[9] ),
    .Y(_07188_));
 inv_2 _11716_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[10] ),
    .Y(_07189_));
 inv_2 _11717_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[11] ),
    .Y(_07190_));
 inv_2 _11718_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[12] ),
    .Y(_07191_));
 inv_2 _11719_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[13] ),
    .Y(_07192_));
 inv_2 _11720_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[14] ),
    .Y(_07193_));
 inv_2 _11721_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[15] ),
    .Y(_07194_));
 inv_2 _11722_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[1] ),
    .Y(_07195_));
 inv_2 _11723_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[1] ),
    .Y(_07196_));
 inv_2 _11724_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[0] ),
    .Y(_07197_));
 inv_2 _11725_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[0] ),
    .Y(_07198_));
 inv_2 _11726_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[2] ),
    .Y(_07199_));
 inv_2 _11727_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[2] ),
    .Y(_07200_));
 inv_2 _11728_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[3] ),
    .Y(_07201_));
 inv_2 _11729_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[3] ),
    .Y(_07202_));
 inv_2 _11730_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[4] ),
    .Y(_07203_));
 inv_2 _11731_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[4] ),
    .Y(_07204_));
 inv_2 _11732_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[5] ),
    .Y(_07205_));
 inv_2 _11733_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[5] ),
    .Y(_07206_));
 inv_2 _11734_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[6] ),
    .Y(_07207_));
 inv_2 _11735_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[6] ),
    .Y(_07208_));
 inv_2 _11736_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key0_r[7] ),
    .Y(_07209_));
 inv_2 _11737_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key1_r[7] ),
    .Y(_07210_));
 inv_2 _11738_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[8] ),
    .Y(_07211_));
 inv_2 _11739_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[9] ),
    .Y(_07212_));
 inv_2 _11740_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[10] ),
    .Y(_07213_));
 inv_2 _11741_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[11] ),
    .Y(_07214_));
 inv_2 _11742_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[12] ),
    .Y(_07215_));
 inv_2 _11743_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[13] ),
    .Y(_07216_));
 inv_2 _11744_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[14] ),
    .Y(_07217_));
 inv_2 _11745_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[15] ),
    .Y(_07218_));
 inv_2 _11746_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[0] ),
    .Y(_07219_));
 inv_2 _11747_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[1] ),
    .Y(_07220_));
 inv_2 _11748_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[2] ),
    .Y(_07221_));
 inv_2 _11749_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[3] ),
    .Y(_07222_));
 inv_2 _11750_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[4] ),
    .Y(_07223_));
 inv_2 _11751_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[5] ),
    .Y(_07224_));
 inv_2 _11752_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[6] ),
    .Y(_07225_));
 inv_2 _11753_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[7] ),
    .Y(_07226_));
 inv_2 _11754_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[0] ),
    .Y(_07227_));
 inv_2 _11755_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[1] ),
    .Y(_07228_));
 inv_2 _11756_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[2] ),
    .Y(_07229_));
 inv_2 _11757_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[3] ),
    .Y(_07230_));
 inv_2 _11758_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[4] ),
    .Y(_07231_));
 inv_2 _11759_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[5] ),
    .Y(_07232_));
 inv_2 _11760_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[6] ),
    .Y(_07233_));
 inv_2 _11761_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key2_r[7] ),
    .Y(_07234_));
 inv_2 _11762_ (.A(\digitop_pav2.sec_inst.shift_in.s9.q[0] ),
    .Y(_07235_));
 inv_2 _11763_ (.A(\digitop_pav2.sync_inst.inst_rstx.gray_counter[2] ),
    .Y(_07236_));
 inv_2 _11764_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m8_clk ),
    .Y(_00158_));
 inv_2 _11765_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m4_clk ),
    .Y(_00157_));
 inv_2 _11766_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m2_clk ),
    .Y(_00156_));
 inv_2 _11767_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.div2 ),
    .Y(_00159_));
 inv_2 _11768_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.div4 ),
    .Y(_00160_));
 inv_2 _11769_ (.A(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.Y ),
    .Y(_00134_));
 inv_2 _11770_ (.A(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.Y ),
    .Y(_00135_));
 inv_2 _11771_ (.A(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.Y ),
    .Y(_00136_));
 inv_2 _11772_ (.A(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.Y ),
    .Y(_00137_));
 inv_2 _11773_ (.A(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.Y ),
    .Y(_00138_));
 inv_2 _11774_ (.A(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.Y ),
    .Y(_00139_));
 inv_2 _11775_ (.A(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.Y ),
    .Y(_00140_));
 inv_2 _11776_ (.A(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.Y ),
    .Y(_00141_));
 inv_2 _11777_ (.A(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.Y ),
    .Y(_00142_));
 inv_2 _11778_ (.A(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.Y ),
    .Y(_00143_));
 inv_2 _11779_ (.A(\digitop_pav2.pie_inst.fsm.clk_i ),
    .Y(_00237_));
 inv_2 _11780_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk4 ),
    .Y(_00132_));
 inv_2 _11781_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk2 ),
    .Y(_00131_));
 inv_2 _11782_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_fc_clk_gated ),
    .Y(_00207_));
 inv_2 _11783_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_en.merge_clk_i ),
    .Y(_00212_));
 inv_2 _11784_ (.A(\digitop_pav2.clkx_irreg_clk ),
    .Y(_00216_));
 inv_2 _11785_ (.A(\digitop_pav2.clkx_invent_clk ),
    .Y(_00248_));
 inv_2 _11786_ (.A(\digitop_pav2.clkx_fm0x_clk ),
    .Y(_00293_));
 inv_2 _11787_ (.A(\digitop_pav2.access_inst.access_ctrl0.nvm_busy_i ),
    .Y(_07237_));
 nor2_1 _11788_ (.A(net1279),
    .B(net1675),
    .Y(_07238_));
 or4_4 _11789_ (.A(net1678),
    .B(net1277),
    .C(net1669),
    .D(net1675),
    .X(_00267_));
 or2_1 _11790_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[5] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state[4] ),
    .X(_07239_));
 nand2_1 _11791_ (.A(_07066_),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state[0] ),
    .Y(_07240_));
 nand2b_2 _11792_ (.A_N(\digitop_pav2.proc_ctrl_inst.cmd.state[3] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state[2] ),
    .Y(_07241_));
 or2_2 _11793_ (.A(_07240_),
    .B(_07241_),
    .X(_07242_));
 nor2_1 _11794_ (.A(net1232),
    .B(_07242_),
    .Y(_07243_));
 or2_4 _11795_ (.A(net1232),
    .B(_07242_),
    .X(_07244_));
 nand2_1 _11796_ (.A(_07065_),
    .B(net1252),
    .Y(_07245_));
 nand2_2 _11797_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[2] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state[3] ),
    .Y(_07246_));
 nor3_1 _11798_ (.A(_07240_),
    .B(net1219),
    .C(_07246_),
    .Y(_07247_));
 or3_4 _11799_ (.A(_07240_),
    .B(net1219),
    .C(_07246_),
    .X(_07248_));
 nor2_1 _11800_ (.A(_07066_),
    .B(net1254),
    .Y(_07249_));
 nand2_1 _11801_ (.A(net1253),
    .B(_07067_),
    .Y(_07250_));
 nor2_1 _11802_ (.A(_07246_),
    .B(_07250_),
    .Y(_07251_));
 and3_2 _11803_ (.A(_07065_),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state[4] ),
    .C(_07251_),
    .X(_07252_));
 nor2_1 _11804_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[2] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state[3] ),
    .Y(_07253_));
 or2_1 _11805_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[2] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state[3] ),
    .X(_07254_));
 nand2_1 _11806_ (.A(_07249_),
    .B(_07253_),
    .Y(_07255_));
 nor2_1 _11807_ (.A(net1219),
    .B(_07255_),
    .Y(_07256_));
 nor2_2 _11808_ (.A(_07252_),
    .B(_07256_),
    .Y(_07257_));
 or2_1 _11809_ (.A(_07252_),
    .B(_07256_),
    .X(_07258_));
 nand2_2 _11810_ (.A(_07248_),
    .B(_07257_),
    .Y(_07259_));
 nand2_4 _11811_ (.A(_07244_),
    .B(_07248_),
    .Y(_07260_));
 nor2_1 _11812_ (.A(net1181),
    .B(_07260_),
    .Y(_07261_));
 nand2_1 _11813_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[5] ),
    .B(net1252),
    .Y(_07262_));
 nand2b_2 _11814_ (.A_N(\digitop_pav2.proc_ctrl_inst.cmd.state[2] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state[3] ),
    .Y(_07263_));
 and4bb_1 _11815_ (.A_N(net1231),
    .B_N(_07263_),
    .C(_07066_),
    .D(_07067_),
    .X(_07264_));
 or4_1 _11816_ (.A(net1253),
    .B(net1254),
    .C(net1231),
    .D(_07263_),
    .X(_07265_));
 nand2_1 _11817_ (.A(net1253),
    .B(net1254),
    .Y(_07266_));
 or2_2 _11818_ (.A(_07246_),
    .B(net1230),
    .X(_07267_));
 inv_2 _11819_ (.A(_07267_),
    .Y(_07268_));
 nor2_1 _11820_ (.A(net1231),
    .B(_07267_),
    .Y(_07269_));
 or2_2 _11821_ (.A(_07264_),
    .B(net1197),
    .X(_07270_));
 or2_1 _11822_ (.A(_07260_),
    .B(_07270_),
    .X(_07271_));
 a21o_1 _11823_ (.A1(net1294),
    .A2(_07271_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdfsm.rn_en ),
    .X(_07272_));
 and2_1 _11824_ (.A(\digitop_pav2.proc_ctrl_inst.inst_checker.state[1] ),
    .B(_07272_),
    .X(_07273_));
 nand2_2 _11825_ (.A(\digitop_pav2.proc_ctrl_inst.inst_checker.state[1] ),
    .B(_07272_),
    .Y(_07274_));
 nor2_1 _11826_ (.A(net1249),
    .B(_07273_),
    .Y(_07275_));
 nand2_2 _11827_ (.A(net1296),
    .B(_07275_),
    .Y(_07276_));
 inv_2 _11828_ (.A(_07276_),
    .Y(_07277_));
 and2_2 _11829_ (.A(net1292),
    .B(_07276_),
    .X(_07278_));
 nand2_1 _11830_ (.A(net1292),
    .B(_07276_),
    .Y(_07279_));
 or4bb_2 _11831_ (.A(net1253),
    .B(net1254),
    .C_N(\digitop_pav2.proc_ctrl_inst.cmd.state[3] ),
    .D_N(\digitop_pav2.proc_ctrl_inst.cmd.state[2] ),
    .X(_07280_));
 nor2_1 _11832_ (.A(net1232),
    .B(_07280_),
    .Y(_07281_));
 or2_1 _11833_ (.A(_07239_),
    .B(_07280_),
    .X(_07282_));
 o21a_2 _11834_ (.A1(net1656),
    .A2(net1251),
    .B1(net1291),
    .X(_07283_));
 and2_1 _11835_ (.A(net1218),
    .B(net1666),
    .X(_07284_));
 nor2_1 _11836_ (.A(net1253),
    .B(_07254_),
    .Y(_07285_));
 nand2_1 _11837_ (.A(_07066_),
    .B(_07253_),
    .Y(_07286_));
 nor2_1 _11838_ (.A(_07065_),
    .B(net1252),
    .Y(_07287_));
 or2_2 _11839_ (.A(_07065_),
    .B(net1252),
    .X(_07288_));
 and3_1 _11840_ (.A(net1254),
    .B(_07285_),
    .C(_07287_),
    .X(_07289_));
 nor2_1 _11841_ (.A(_07270_),
    .B(net1196),
    .Y(_07290_));
 or2_1 _11842_ (.A(_07270_),
    .B(net1196),
    .X(_07291_));
 nor2_4 _11843_ (.A(_07267_),
    .B(_07288_),
    .Y(_07292_));
 or2_2 _11844_ (.A(_07267_),
    .B(_07288_),
    .X(_07293_));
 nor2_1 _11845_ (.A(net1181),
    .B(_07292_),
    .Y(_07294_));
 nand2_2 _11846_ (.A(_07257_),
    .B(_07293_),
    .Y(_07295_));
 or3_2 _11847_ (.A(_07247_),
    .B(_07291_),
    .C(_07295_),
    .X(_07296_));
 nand2_1 _11848_ (.A(net1291),
    .B(_07296_),
    .Y(_07297_));
 and2_2 _11849_ (.A(net1666),
    .B(_07296_),
    .X(_07298_));
 nor2_2 _11850_ (.A(_07284_),
    .B(_07298_),
    .Y(_07299_));
 or3_1 _11851_ (.A(_07256_),
    .B(_07264_),
    .C(net1196),
    .X(_07300_));
 or2_1 _11852_ (.A(_07256_),
    .B(_07291_),
    .X(_07301_));
 or2_1 _11853_ (.A(net1186),
    .B(_07252_),
    .X(_07302_));
 or2_1 _11854_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[0] ),
    .B(_07241_),
    .X(_07303_));
 or2_1 _11855_ (.A(net1253),
    .B(_07303_),
    .X(_07304_));
 nor2_1 _11856_ (.A(net1219),
    .B(_07304_),
    .Y(_07305_));
 inv_2 _11857_ (.A(net1185),
    .Y(_07306_));
 nand2_1 _11858_ (.A(net1254),
    .B(_07253_),
    .Y(_07307_));
 nor2_1 _11859_ (.A(_07254_),
    .B(net1230),
    .Y(_07308_));
 or2_1 _11860_ (.A(_07254_),
    .B(net1230),
    .X(_07309_));
 nor2_2 _11861_ (.A(_07239_),
    .B(_07309_),
    .Y(_07310_));
 or2_2 _11862_ (.A(net1232),
    .B(_07309_),
    .X(_07311_));
 nor2_1 _11863_ (.A(net1185),
    .B(net1195),
    .Y(_07312_));
 or2_2 _11864_ (.A(net1185),
    .B(_07310_),
    .X(_07313_));
 or3_1 _11865_ (.A(net1198),
    .B(_07292_),
    .C(_07313_),
    .X(_07314_));
 or2_1 _11866_ (.A(_07302_),
    .B(_07314_),
    .X(_07315_));
 or2_1 _11867_ (.A(_07301_),
    .B(_07315_),
    .X(_07316_));
 and2_1 _11868_ (.A(net1288),
    .B(_07252_),
    .X(_07317_));
 and2_1 _11869_ (.A(net1288),
    .B(_07314_),
    .X(_07318_));
 nand2_1 _11870_ (.A(net1286),
    .B(_07316_),
    .Y(_07319_));
 nor2_1 _11871_ (.A(net1262),
    .B(net1699),
    .Y(_07320_));
 or2_1 _11872_ (.A(net1260),
    .B(net1699),
    .X(_07321_));
 and3_1 _11873_ (.A(net1239),
    .B(net1695),
    .C(_07320_),
    .X(_07322_));
 inv_2 _11874_ (.A(net1211),
    .Y(\digitop_pav2.sync_inst.inst_clkx.g_access ));
 or2_2 _11875_ (.A(net1691),
    .B(_00267_),
    .X(_00168_));
 or2_1 _11876_ (.A(net1626),
    .B(net1658),
    .X(_07323_));
 nor4_1 _11877_ (.A(net1273),
    .B(_00267_),
    .C(net1194),
    .D(_07323_),
    .Y(_07324_));
 or3_2 _11878_ (.A(\digitop_pav2.sync_inst.inst_clkx.g_access ),
    .B(net1199),
    .C(_07323_),
    .X(_07325_));
 o211a_1 _11879_ (.A1(net1198),
    .A2(net1659),
    .B1(_07260_),
    .C1(net1294),
    .X(_07326_));
 or2_2 _11880_ (.A(net1643),
    .B(net1721),
    .X(_07327_));
 nor2_2 _11881_ (.A(_07087_),
    .B(net1215),
    .Y(_07328_));
 nand2_1 _11882_ (.A(net1286),
    .B(net1217),
    .Y(_07329_));
 nor2_1 _11883_ (.A(net1218),
    .B(_07313_),
    .Y(_07330_));
 nand2_1 _11884_ (.A(net1215),
    .B(_07312_),
    .Y(_07331_));
 nor2_1 _11885_ (.A(net1218),
    .B(_07314_),
    .Y(_07332_));
 o211a_1 _11886_ (.A1(_07261_),
    .A2(net1663),
    .B1(_07319_),
    .C1(_07329_),
    .X(_07333_));
 and4bb_4 _11887_ (.A_N(net1660),
    .B_N(net1644),
    .C(net1664),
    .D(_07299_),
    .X(_07334_));
 or4bb_1 _11888_ (.A(net1660),
    .B(net1644),
    .C_N(_07333_),
    .D_N(_07299_),
    .X(_07335_));
 and3_2 _11889_ (.A(net1248),
    .B(_00267_),
    .C(net818),
    .X(_07336_));
 or3b_1 _11890_ (.A(_07334_),
    .B(net1233),
    .C_N(_00267_),
    .X(_07337_));
 nor2_1 _11891_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[9] ),
    .B(net1172),
    .Y(_07338_));
 or2_4 _11892_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[9] ),
    .B(net1172),
    .X(_07339_));
 mux2_1 _11893_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[3] ),
    .A1(_07339_),
    .S(_07336_),
    .X(_01605_));
 mux2_1 _11894_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[6] ),
    .A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[5] ),
    .S(net808),
    .X(_01604_));
 mux2_1 _11895_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[13] ),
    .A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[9] ),
    .S(net808),
    .X(_01603_));
 mux2_1 _11896_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[13] ),
    .A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[11] ),
    .S(_07336_),
    .X(_01602_));
 or3_1 _11897_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[6] ),
    .B(\digitop_pav2.access_inst.access_check0.wordcnt_i[4] ),
    .C(\digitop_pav2.access_inst.access_check0.wordcnt_i[5] ),
    .X(_07340_));
 nor4_1 _11898_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[1] ),
    .B(\digitop_pav2.access_inst.access_check0.wordcnt_i[2] ),
    .C(\digitop_pav2.access_inst.access_check0.wordcnt_i[3] ),
    .D(_07340_),
    .Y(_07341_));
 nor2_1 _11899_ (.A(_07038_),
    .B(net1238),
    .Y(_07342_));
 o21a_1 _11900_ (.A1(\digitop_pav2.access_inst.access_ctrl0.state[25] ),
    .A2(net1143),
    .B1(_07342_),
    .X(_07343_));
 o21ai_2 _11901_ (.A1(\digitop_pav2.access_inst.access_ctrl0.state[25] ),
    .A2(net1143),
    .B1(_07342_),
    .Y(_07344_));
 o21ai_1 _11902_ (.A1(net1071),
    .A2(\digitop_pav2.access_inst.access_check0.wordcnt_i[0] ),
    .B1(net1650),
    .Y(_07345_));
 a21oi_1 _11903_ (.A1(net1071),
    .A2(\digitop_pav2.access_inst.access_check0.wordcnt_i[0] ),
    .B1(_07345_),
    .Y(_07346_));
 a31o_1 _11904_ (.A1(net1018),
    .A2(net1011),
    .A3(_07346_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.proc_rd_finish_i ),
    .X(_01584_));
 and2_1 _11905_ (.A(net1303),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[11] ),
    .X(_07347_));
 and2_1 _11906_ (.A(net1303),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[4] ),
    .X(_07348_));
 nor2_1 _11907_ (.A(net1710),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[4] ),
    .Y(_07349_));
 or2_1 _11908_ (.A(net1710),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[4] ),
    .X(_07350_));
 and2_1 _11909_ (.A(net1304),
    .B(net1290),
    .X(_07351_));
 nand2_4 _11910_ (.A(net1304),
    .B(net1290),
    .Y(_07352_));
 or3_1 _11911_ (.A(_07291_),
    .B(_07295_),
    .C(_07331_),
    .X(_07353_));
 nor2_1 _11912_ (.A(_07290_),
    .B(_07352_),
    .Y(_07354_));
 a22o_1 _11913_ (.A1(net1303),
    .A2(_07350_),
    .B1(net1229),
    .B2(_07353_),
    .X(_07355_));
 or4_1 _11914_ (.A(\digitop_pav2.proc_ctrl_inst.ebv.state[4] ),
    .B(\digitop_pav2.proc_ctrl_inst.ebv.state[2] ),
    .C(\digitop_pav2.proc_ctrl_inst.ebv.state[9] ),
    .D(\digitop_pav2.proc_ctrl_inst.ebv.state[5] ),
    .X(_07356_));
 or4_1 _11915_ (.A(\digitop_pav2.proc_ctrl_inst.ebv.state[12] ),
    .B(\digitop_pav2.proc_ctrl_inst.ebv.state[10] ),
    .C(\digitop_pav2.proc_ctrl_inst.ebv.state[14] ),
    .D(_07356_),
    .X(_07357_));
 and2_1 _11916_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[4] ),
    .B(net971),
    .X(_07358_));
 a221o_1 _11917_ (.A1(net1710),
    .A2(_07295_),
    .B1(_07357_),
    .B2(_07358_),
    .C1(_07349_),
    .X(_07359_));
 or3_2 _11918_ (.A(net1218),
    .B(net1196),
    .C(net1185),
    .X(_07360_));
 nand2_2 _11919_ (.A(net1215),
    .B(_07293_),
    .Y(_07361_));
 or3_1 _11920_ (.A(_07295_),
    .B(net1195),
    .C(_07360_),
    .X(_07362_));
 o41a_4 _11921_ (.A1(net1273),
    .A2(_00267_),
    .A3(\digitop_pav2.sync_inst.inst_clkx.g_access ),
    .A4(_07323_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[0] ),
    .X(_07363_));
 nand2_1 _11922_ (.A(_07257_),
    .B(net1184),
    .Y(_07364_));
 and4_1 _11923_ (.A(net1216),
    .B(_07293_),
    .C(_07311_),
    .D(_07363_),
    .X(_07365_));
 o31a_1 _11924_ (.A1(net1196),
    .A2(_07313_),
    .A3(_07361_),
    .B1(_07363_),
    .X(_07366_));
 and3_1 _11925_ (.A(net1295),
    .B(_07362_),
    .C(_07364_),
    .X(_07367_));
 a22oi_4 _11926_ (.A1(_07355_),
    .A2(net1711),
    .B1(_07367_),
    .B2(net1303),
    .Y(_07368_));
 a21oi_1 _11927_ (.A1(\digitop_pav2.access_inst.access_ctrl0.rx_par0_i ),
    .A2(net1702),
    .B1(\digitop_pav2.access_inst.access_ctrl0.state[17] ),
    .Y(_07369_));
 nor2_1 _11928_ (.A(net1712),
    .B(_07369_),
    .Y(_07370_));
 o21a_1 _11929_ (.A1(\digitop_pav2.access_inst.access_ctrl0.state[13] ),
    .A2(\digitop_pav2.access_inst.access_ctrl0.state[17] ),
    .B1(_07370_),
    .X(_07371_));
 or2_2 _11930_ (.A(\digitop_pav2.access_inst.access_check0.mem_sign_check_i ),
    .B(\digitop_pav2.access_inst.access_check0.pc_lock_check_i ),
    .X(_07372_));
 nor2_2 _11931_ (.A(net1210),
    .B(_07372_),
    .Y(_07373_));
 and2b_1 _11932_ (.A_N(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[1] ),
    .B(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[0] ),
    .X(_07374_));
 and2b_2 _11933_ (.A_N(net1042),
    .B(net1040),
    .X(_07375_));
 and2_2 _11934_ (.A(_07374_),
    .B(_07375_),
    .X(_07376_));
 a31o_1 _11935_ (.A1(_07371_),
    .A2(_07373_),
    .A3(_07376_),
    .B1(\digitop_pav2.access_inst.access_transceiver0.wcnt_stb_valid ),
    .X(_01567_));
 a31o_1 _11936_ (.A1(_07349_),
    .A2(net1229),
    .A3(_07353_),
    .B1(_07367_),
    .X(_07377_));
 and3_1 _11937_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[11] ),
    .B(net1638),
    .C(_07295_),
    .X(_07378_));
 o22a_1 _11938_ (.A1(net1638),
    .A2(\digitop_pav2.proc_ctrl_inst.ebv.invalid ),
    .B1(_07358_),
    .B2(_07378_),
    .X(_07379_));
 a32o_1 _11939_ (.A1(net1303),
    .A2(_07350_),
    .A3(_07379_),
    .B1(_07377_),
    .B2(net1638),
    .X(_07380_));
 a41o_1 _11940_ (.A1(net1702),
    .A2(_07370_),
    .A3(_07376_),
    .A4(net1640),
    .B1(\digitop_pav2.access_inst.access_check0.error_wordcnt_i ),
    .X(_01566_));
 and3_1 _11941_ (.A(\digitop_pav2.access_inst.access_ctrl0.replay_ok ),
    .B(net1702),
    .C(net1142),
    .X(_07381_));
 a21oi_1 _11942_ (.A1(\digitop_pav2.access_inst.access_ctrl0.replay_nok ),
    .A2(net1142),
    .B1(_07381_),
    .Y(_07382_));
 and2_1 _11943_ (.A(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[1] ),
    .B(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[0] ),
    .X(_07383_));
 and3_1 _11944_ (.A(net1042),
    .B(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[1] ),
    .C(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[0] ),
    .X(_07384_));
 and2_1 _11945_ (.A(net1040),
    .B(_07384_),
    .X(_07385_));
 nand2_1 _11946_ (.A(net1041),
    .B(_07384_),
    .Y(_07386_));
 or4_2 _11947_ (.A(\digitop_pav2.access_inst.access_ctrl0.state[15] ),
    .B(net1142),
    .C(net1143),
    .D(\digitop_pav2.access_inst.access_ctrl0.state[22] ),
    .X(_07387_));
 a41o_1 _11948_ (.A1(_07373_),
    .A2(_07382_),
    .A3(_07385_),
    .A4(_07387_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.dt_acc_done_o ),
    .X(_01565_));
 and3_1 _11949_ (.A(\digitop_pav2.access_inst.access_ctrl0.replay_nok ),
    .B(net1142),
    .C(_07384_),
    .X(_07388_));
 nand2_2 _11950_ (.A(_07053_),
    .B(net1018),
    .Y(_07389_));
 nor2_1 _11951_ (.A(_07386_),
    .B(_07389_),
    .Y(_07390_));
 a31o_1 _11952_ (.A1(\digitop_pav2.access_inst.access_ctrl0.proc_rd_finish_i ),
    .A2(_07381_),
    .A3(_07390_),
    .B1(_07388_),
    .X(_07391_));
 a21o_1 _11953_ (.A1(_07373_),
    .A2(_07391_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.tx_dt_finish_i ),
    .X(_01548_));
 nor2_1 _11954_ (.A(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[1] ),
    .B(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[0] ),
    .Y(_07392_));
 nor2_2 _11955_ (.A(net1040),
    .B(net1042),
    .Y(_07393_));
 and2_1 _11956_ (.A(_07392_),
    .B(_07393_),
    .X(_07394_));
 a31o_1 _11957_ (.A1(_07371_),
    .A2(_07373_),
    .A3(_07394_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.rx_par1_i ),
    .X(_01547_));
 nor2_2 _11958_ (.A(net1699),
    .B(net1694),
    .Y(_07395_));
 or2_2 _11959_ (.A(net1699),
    .B(net1694),
    .X(_07396_));
 o21a_1 _11960_ (.A1(net1702),
    .A2(_07396_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.state[0] ),
    .X(_07397_));
 nand2_1 _11961_ (.A(\digitop_pav2.access_inst.access_ctrl0.rx_par0_i ),
    .B(_07396_),
    .Y(_07398_));
 a21oi_1 _11962_ (.A1(\digitop_pav2.access_inst.access_ctrl0.state[13] ),
    .A2(_07398_),
    .B1(_07397_),
    .Y(_07399_));
 nor2_1 _11963_ (.A(net1712),
    .B(_07399_),
    .Y(_07400_));
 or4_1 _11964_ (.A(\digitop_pav2.access_inst.access_ctrl0.state[13] ),
    .B(\digitop_pav2.access_inst.access_ctrl0.state[20] ),
    .C(\digitop_pav2.access_inst.access_ctrl0.state[17] ),
    .D(_07397_),
    .X(_07401_));
 nand2_1 _11965_ (.A(_07375_),
    .B(_07392_),
    .Y(_07402_));
 o21a_1 _11966_ (.A1(\digitop_pav2.access_inst.access_ctrl0.state[13] ),
    .A2(\digitop_pav2.access_inst.access_ctrl0.state[0] ),
    .B1(net1694),
    .X(_07403_));
 nor2_1 _11967_ (.A(_07402_),
    .B(_07403_),
    .Y(_07404_));
 and2b_2 _11968_ (.A_N(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[0] ),
    .B(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[1] ),
    .X(_07405_));
 and3b_1 _11969_ (.A_N(net1040),
    .B(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[2] ),
    .C(_07405_),
    .X(_07406_));
 a21o_1 _11970_ (.A1(_07403_),
    .A2(_07406_),
    .B1(_07404_),
    .X(_07407_));
 a41o_1 _11971_ (.A1(_07373_),
    .A2(_07400_),
    .A3(_07401_),
    .A4(_07407_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.rx_par0_i ),
    .X(_01546_));
 o21a_1 _11972_ (.A1(_07395_),
    .A2(_07399_),
    .B1(net1194),
    .X(_07408_));
 and3_1 _11973_ (.A(_07334_),
    .B(_07387_),
    .C(_07408_),
    .X(_07409_));
 or2_1 _11974_ (.A(\digitop_pav2.access_inst.access_ctrl0.state[15] ),
    .B(net1142),
    .X(_07410_));
 or2_1 _11975_ (.A(\digitop_pav2.access_inst.access_ctrl0.tx_dt_finish_i ),
    .B(_07382_),
    .X(_07411_));
 nand2_1 _11976_ (.A(_07410_),
    .B(_07411_),
    .Y(_07412_));
 o21a_1 _11977_ (.A1(net1042),
    .A2(_07090_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.replay_nok ),
    .X(_07413_));
 mux2_1 _11978_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[15] ),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[15] ),
    .S(net1045),
    .X(_07414_));
 and3_1 _11979_ (.A(net1040),
    .B(net1042),
    .C(_07392_),
    .X(_07415_));
 and3b_1 _11980_ (.A_N(net1040),
    .B(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[2] ),
    .C(_07374_),
    .X(_07416_));
 mux2_1 _11981_ (.A0(\digitop_pav2.boot_inst.boot_proc0.proc_fg[12] ),
    .A1(_07100_),
    .S(\digitop_pav2.access_inst.access_check0.fg_i[8] ),
    .X(_07417_));
 mux2_1 _11982_ (.A0(_07101_),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[3] ),
    .S(\digitop_pav2.access_inst.access_check0.fg_i[8] ),
    .X(_07418_));
 and3_1 _11983_ (.A(_07393_),
    .B(_07405_),
    .C(net1318),
    .X(_07419_));
 and2b_1 _11984_ (.A_N(net1040),
    .B(_07384_),
    .X(_07420_));
 and3_1 _11985_ (.A(net1040),
    .B(net1042),
    .C(_07405_),
    .X(_07421_));
 and3_1 _11986_ (.A(net1040),
    .B(net1042),
    .C(_07374_),
    .X(_07422_));
 and3b_1 _11987_ (.A_N(net1040),
    .B(net1042),
    .C(_07392_),
    .X(_07423_));
 a22o_1 _11988_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[1] ),
    .A2(_07422_),
    .B1(_07423_),
    .B2(\digitop_pav2.access_inst.access_check0.fg_i[10] ),
    .X(_07424_));
 a2bb2o_1 _11989_ (.A1_N(_07098_),
    .A2_N(_07402_),
    .B1(_07415_),
    .B2(\digitop_pav2.access_inst.access_check0.fg_i[2] ),
    .X(_07425_));
 a32o_1 _11990_ (.A1(net1323),
    .A2(_07375_),
    .A3(_07405_),
    .B1(_07420_),
    .B2(\digitop_pav2.access_inst.access_check0.fg_i[7] ),
    .X(_07426_));
 a311o_1 _11991_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[3] ),
    .A2(_07375_),
    .A3(_07383_),
    .B1(_07419_),
    .C1(_07426_),
    .X(_07427_));
 a221o_1 _11992_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[8] ),
    .A2(_07406_),
    .B1(_07421_),
    .B2(\digitop_pav2.access_inst.access_check0.fg_i[0] ),
    .C1(_07424_),
    .X(_07428_));
 a221o_1 _11993_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[5] ),
    .A2(_07376_),
    .B1(_07416_),
    .B2(\digitop_pav2.access_inst.access_check0.fg_i[9] ),
    .C1(_07428_),
    .X(_07429_));
 a311o_1 _11994_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[11] ),
    .A2(_07383_),
    .A3(_07393_),
    .B1(_07427_),
    .C1(_07429_),
    .X(_07430_));
 a31o_1 _11995_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[13] ),
    .A2(_07374_),
    .A3(_07393_),
    .B1(net1695),
    .X(_07431_));
 a32o_1 _11996_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[14] ),
    .A2(_07374_),
    .A3(_07393_),
    .B1(_07376_),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[6] ),
    .X(_07432_));
 and3_1 _11997_ (.A(\digitop_pav2.access_inst.access_transceiver0.handle_i[4] ),
    .B(_07375_),
    .C(_07383_),
    .X(_07433_));
 a311o_1 _11998_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[13] ),
    .A2(_07393_),
    .A3(_07405_),
    .B1(_07432_),
    .C1(_07433_),
    .X(_07434_));
 a22o_1 _11999_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[10] ),
    .A2(_07416_),
    .B1(_07422_),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[2] ),
    .X(_07435_));
 a21o_1 _12000_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[8] ),
    .A2(_07420_),
    .B1(_07435_),
    .X(_07436_));
 a32o_1 _12001_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[5] ),
    .A2(_07375_),
    .A3(_07405_),
    .B1(_07385_),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[0] ),
    .X(_07437_));
 a221o_1 _12002_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[9] ),
    .A2(_07406_),
    .B1(_07415_),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[3] ),
    .C1(_07437_),
    .X(_07438_));
 and3_1 _12003_ (.A(\digitop_pav2.access_inst.access_transceiver0.handle_i[7] ),
    .B(_07375_),
    .C(_07392_),
    .X(_07439_));
 a31o_1 _12004_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[12] ),
    .A2(_07383_),
    .A3(_07393_),
    .B1(_07439_),
    .X(_07440_));
 a221o_1 _12005_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[1] ),
    .A2(_07421_),
    .B1(_07423_),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[11] ),
    .C1(_07440_),
    .X(_07441_));
 or4_1 _12006_ (.A(_07434_),
    .B(_07436_),
    .C(_07438_),
    .D(_07441_),
    .X(_07442_));
 a211o_1 _12007_ (.A1(net1729),
    .A2(_07394_),
    .B1(_07442_),
    .C1(net1694),
    .X(_07443_));
 o31a_1 _12008_ (.A1(_07425_),
    .A2(_07430_),
    .A3(_07431_),
    .B1(net1730),
    .X(_07444_));
 mux2_1 _12009_ (.A0(_07413_),
    .A1(_07414_),
    .S(_07381_),
    .X(_07445_));
 o311a_1 _12010_ (.A1(net1240),
    .A2(net1142),
    .A3(\digitop_pav2.access_inst.access_ctrl0.state[22] ),
    .B1(_07412_),
    .C1(_07445_),
    .X(_07446_));
 a31o_1 _12011_ (.A1(_07410_),
    .A2(_07411_),
    .A3(net1731),
    .B1(_07446_),
    .X(_07447_));
 mux2_1 _12012_ (.A0(\digitop_pav2.access_inst.access_ctrl0.tx_bit_i ),
    .A1(_07447_),
    .S(_07409_),
    .X(_01545_));
 nor2_1 _12013_ (.A(net1194),
    .B(_07372_),
    .Y(_07448_));
 a31o_1 _12014_ (.A1(\digitop_pav2.access_inst.access_ctrl0.rx_par0_i ),
    .A2(\digitop_pav2.access_inst.access_ctrl0.state[13] ),
    .A3(_07396_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.state[20] ),
    .X(_07449_));
 and2b_1 _12015_ (.A_N(net1712),
    .B(_07449_),
    .X(_07450_));
 a31o_1 _12016_ (.A1(net1276),
    .A2(_07334_),
    .A3(_07450_),
    .B1(_07371_),
    .X(_07451_));
 nand2_1 _12017_ (.A(net1699),
    .B(_07404_),
    .Y(_07452_));
 nor2_1 _12018_ (.A(_07400_),
    .B(_07451_),
    .Y(_07453_));
 a21o_1 _12019_ (.A1(_07400_),
    .A2(_07452_),
    .B1(_07451_),
    .X(_07454_));
 xor2_1 _12020_ (.A(net1041),
    .B(_07384_),
    .X(_07455_));
 o31a_1 _12021_ (.A1(_07037_),
    .A2(_07090_),
    .A3(_07342_),
    .B1(_07387_),
    .X(_07456_));
 a22o_1 _12022_ (.A1(net1041),
    .A2(_07453_),
    .B1(_07454_),
    .B2(_07455_),
    .X(_07457_));
 nand2_1 _12023_ (.A(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[0] ),
    .B(_07410_),
    .Y(_07458_));
 nand2_1 _12024_ (.A(_07384_),
    .B(_07410_),
    .Y(_07459_));
 xnor2_1 _12025_ (.A(net1041),
    .B(_07459_),
    .Y(_07460_));
 mux2_1 _12026_ (.A0(_07457_),
    .A1(_07460_),
    .S(_07456_),
    .X(_07461_));
 a22o_1 _12027_ (.A1(net1041),
    .A2(_07448_),
    .B1(_07461_),
    .B2(_07373_),
    .X(_01544_));
 o21a_1 _12028_ (.A1(_07400_),
    .A2(_07451_),
    .B1(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[0] ),
    .X(_07462_));
 inv_2 _12029_ (.A(_07462_),
    .Y(_07463_));
 nand2_1 _12030_ (.A(_07387_),
    .B(_07458_),
    .Y(_07464_));
 o211a_1 _12031_ (.A1(_07387_),
    .A2(_07462_),
    .B1(_07464_),
    .C1(net1194),
    .X(_07465_));
 and2_1 _12032_ (.A(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[1] ),
    .B(_07465_),
    .X(_07466_));
 a31o_1 _12033_ (.A1(net1042),
    .A2(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[1] ),
    .A3(_07465_),
    .B1(_07372_),
    .X(_07467_));
 o21ba_1 _12034_ (.A1(net1042),
    .A2(_07466_),
    .B1_N(_07467_),
    .X(_01543_));
 nor2_1 _12035_ (.A(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[1] ),
    .B(_07465_),
    .Y(_07468_));
 nor3_1 _12036_ (.A(_07372_),
    .B(_07466_),
    .C(_07468_),
    .Y(_01542_));
 or2_1 _12037_ (.A(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[0] ),
    .B(_07454_),
    .X(_07469_));
 a21o_1 _12038_ (.A1(_07463_),
    .A2(_07469_),
    .B1(_07387_),
    .X(_07470_));
 or2_1 _12039_ (.A(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[0] ),
    .B(_07410_),
    .X(_07471_));
 a21bo_1 _12040_ (.A1(_07458_),
    .A2(_07471_),
    .B1_N(_07387_),
    .X(_07472_));
 a32o_1 _12041_ (.A1(_07373_),
    .A2(_07470_),
    .A3(_07472_),
    .B1(_07448_),
    .B2(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[0] ),
    .X(_01541_));
 nand2_1 _12042_ (.A(_07373_),
    .B(_07381_),
    .Y(_07473_));
 nor2_1 _12043_ (.A(_07386_),
    .B(_07473_),
    .Y(_07474_));
 xor2_1 _12044_ (.A(net1045),
    .B(_07474_),
    .X(_01540_));
 mux2_1 _12045_ (.A0(_07394_),
    .A1(\digitop_pav2.access_inst.access_ctrl0.tx_proc_rd_stb_i ),
    .S(_07473_),
    .X(_01539_));
 nor2_1 _12046_ (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[1] ),
    .B(net1049),
    .Y(_07475_));
 or2_2 _12047_ (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[1] ),
    .B(net1049),
    .X(_07476_));
 nor2_4 _12048_ (.A(net1155),
    .B(_07476_),
    .Y(_07477_));
 nand2_1 _12049_ (.A(net1036),
    .B(_07475_),
    .Y(_07478_));
 nand2_2 _12050_ (.A(_07031_),
    .B(_07477_),
    .Y(_07479_));
 nor2_2 _12051_ (.A(net1240),
    .B(net1235),
    .Y(_07480_));
 nand2_1 _12052_ (.A(net1258),
    .B(net1650),
    .Y(_07481_));
 nor3_1 _12053_ (.A(\digitop_pav2.access_inst.access_ctrl0.state[9] ),
    .B(\digitop_pav2.access_inst.access_ctrl0.state[2] ),
    .C(\digitop_pav2.access_inst.access_check0.wr_lock_ck_i ),
    .Y(_07482_));
 or3_2 _12054_ (.A(\digitop_pav2.access_inst.access_ctrl0.state[9] ),
    .B(\digitop_pav2.access_inst.access_ctrl0.state[2] ),
    .C(\digitop_pav2.access_inst.access_check0.wr_lock_ck_i ),
    .X(_07483_));
 or4_1 _12055_ (.A(net1148),
    .B(net1152),
    .C(\digitop_pav2.access_inst.access_ctrl0.state[11] ),
    .D(\digitop_pav2.access_inst.access_ctrl0.state[10] ),
    .X(_07484_));
 or4_1 _12056_ (.A(net1144),
    .B(net1145),
    .C(\digitop_pav2.access_inst.access_ctrl0.state[23] ),
    .D(_07484_),
    .X(_07485_));
 or4_1 _12057_ (.A(\digitop_pav2.access_inst.access_ctrl0.state[24] ),
    .B(\digitop_pav2.access_inst.access_ctrl0.state[14] ),
    .C(\digitop_pav2.access_inst.access_ctrl0.ld_dt_stb ),
    .D(\digitop_pav2.access_inst.access_ctrl0.state[18] ),
    .X(_07486_));
 nor4_1 _12058_ (.A(net1011),
    .B(_07483_),
    .C(_07485_),
    .D(_07486_),
    .Y(_07487_));
 or4_4 _12059_ (.A(net1011),
    .B(_07483_),
    .C(_07485_),
    .D(_07486_),
    .X(_07488_));
 or3_2 _12060_ (.A(_07481_),
    .B(_07483_),
    .C(net964),
    .X(_07489_));
 nor2_1 _12061_ (.A(_07479_),
    .B(_07489_),
    .Y(_07490_));
 nor2_2 _12062_ (.A(_07024_),
    .B(net1065),
    .Y(_07491_));
 nand2_1 _12063_ (.A(_07030_),
    .B(net1065),
    .Y(_07492_));
 nor2_2 _12064_ (.A(\digitop_pav2.access_inst.access_check0.ctrl_wcknzero_ck ),
    .B(_07492_),
    .Y(_07493_));
 nand2_1 _12065_ (.A(net1046),
    .B(net1258),
    .Y(_07494_));
 nor3_1 _12066_ (.A(_07491_),
    .B(_07493_),
    .C(_07494_),
    .Y(_07495_));
 a31o_1 _12067_ (.A1(net1063),
    .A2(_07490_),
    .A3(_07495_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.ld_key_env_finish_i ),
    .X(_01538_));
 nor2_1 _12068_ (.A(\digitop_pav2.access_inst.access_ctrl0.nvm_busy_i ),
    .B(_07476_),
    .Y(_07496_));
 a41o_1 _12069_ (.A1(_07480_),
    .A2(_07482_),
    .A3(net963),
    .A4(_07496_),
    .B1(net1047),
    .X(_01537_));
 nor2_4 _12070_ (.A(net1239),
    .B(net1034),
    .Y(_07497_));
 nand2_2 _12071_ (.A(net1257),
    .B(_07483_),
    .Y(_07498_));
 nand2_1 _12072_ (.A(_07069_),
    .B(_07498_),
    .Y(_07499_));
 o211a_1 _12073_ (.A1(net1047),
    .A2(net1063),
    .B1(net1065),
    .C1(net1257),
    .X(_07500_));
 and4_1 _12074_ (.A(_07023_),
    .B(_07033_),
    .C(net1069),
    .D(_07500_),
    .X(_07501_));
 a21o_1 _12075_ (.A1(net1239),
    .A2(\digitop_pav2.access_inst.access_transceiver0.rx_par_buf[15] ),
    .B1(_07501_),
    .X(_07502_));
 nor2_4 _12076_ (.A(_07499_),
    .B(_07502_),
    .Y(_07503_));
 or2_2 _12077_ (.A(_07499_),
    .B(_07502_),
    .X(_07504_));
 a21o_1 _12078_ (.A1(net1047),
    .A2(\digitop_pav2.access_inst.access_ctrl0.crc_init_i ),
    .B1(net1239),
    .X(_07505_));
 nand2_1 _12079_ (.A(net1239),
    .B(\digitop_pav2.access_inst.access_transceiver0.rx_par_buf[14] ),
    .Y(_07506_));
 o22a_1 _12080_ (.A1(net1069),
    .A2(net1239),
    .B1(_07505_),
    .B2(net1065),
    .X(_07507_));
 a21o_1 _12081_ (.A1(_07506_),
    .A2(_07507_),
    .B1(_07499_),
    .X(_07508_));
 inv_2 _12082_ (.A(net962),
    .Y(_07509_));
 nor2_4 _12083_ (.A(_07503_),
    .B(_07509_),
    .Y(_07510_));
 nand2_4 _12084_ (.A(_07504_),
    .B(net962),
    .Y(_07511_));
 and2_1 _12085_ (.A(net1156),
    .B(net1157),
    .X(_07512_));
 nand2_2 _12086_ (.A(net1156),
    .B(net1157),
    .Y(_07513_));
 or2_1 _12087_ (.A(net1156),
    .B(net1157),
    .X(_07514_));
 and4_1 _12088_ (.A(_07031_),
    .B(net1260),
    .C(_07513_),
    .D(_07514_),
    .X(_07515_));
 nor2_1 _12089_ (.A(net471),
    .B(net431),
    .Y(_07516_));
 or2_4 _12090_ (.A(net473),
    .B(net439),
    .X(_07517_));
 or2_1 _12091_ (.A(net470),
    .B(net426),
    .X(_07518_));
 nor2_1 _12092_ (.A(_07517_),
    .B(_07518_),
    .Y(_07519_));
 or2_4 _12093_ (.A(_07517_),
    .B(_07518_),
    .X(_07520_));
 or3_1 _12094_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[4] ),
    .C(net463),
    .X(_07521_));
 nor2_1 _12095_ (.A(_07520_),
    .B(_07521_),
    .Y(_07522_));
 or2_2 _12096_ (.A(_07520_),
    .B(_07521_),
    .X(_07523_));
 nor2_2 _12097_ (.A(_07023_),
    .B(_07523_),
    .Y(_07524_));
 nand2_1 _12098_ (.A(net1256),
    .B(_07524_),
    .Y(_07525_));
 o211a_1 _12099_ (.A1(net1066),
    .A2(_07525_),
    .B1(_07515_),
    .C1(net962),
    .X(_07526_));
 nor2_1 _12100_ (.A(_07504_),
    .B(net962),
    .Y(_07527_));
 or2_2 _12101_ (.A(_07504_),
    .B(net962),
    .X(_07528_));
 nor2_1 _12102_ (.A(net1073),
    .B(net1074),
    .Y(_07529_));
 or2_1 _12103_ (.A(\digitop_pav2.access_inst.access_check0.wordptr_i[5] ),
    .B(net1074),
    .X(_07530_));
 nor2_1 _12104_ (.A(net1072),
    .B(_07530_),
    .Y(_07531_));
 or2_1 _12105_ (.A(net1072),
    .B(_07530_),
    .X(_07532_));
 nor2_1 _12106_ (.A(net1081),
    .B(net1079),
    .Y(_07533_));
 nor2_1 _12107_ (.A(net1077),
    .B(net1075),
    .Y(_07534_));
 nor2_1 _12108_ (.A(net1079),
    .B(net1077),
    .Y(_07535_));
 or3_1 _12109_ (.A(net1081),
    .B(net1079),
    .C(net1077),
    .X(_07536_));
 or2_1 _12110_ (.A(net1075),
    .B(_07536_),
    .X(_07537_));
 nor2_1 _12111_ (.A(_07532_),
    .B(_07537_),
    .Y(_07538_));
 or2_1 _12112_ (.A(_07532_),
    .B(_07537_),
    .X(_07539_));
 o2111a_1 _12113_ (.A1(\digitop_pav2.access_inst.access_check0.wcnt_check_zero ),
    .A2(net1037),
    .B1(net913),
    .C1(_07538_),
    .D1(\digitop_pav2.access_inst.access_ctrl0.tx_proc_rd_stb_i ),
    .X(_07540_));
 a211oi_1 _12114_ (.A1(net1037),
    .A2(_07540_),
    .B1(_07536_),
    .C1(net1257),
    .Y(_07541_));
 or3b_1 _12115_ (.A(net1056),
    .B(net1058),
    .C_N(net1060),
    .X(_07542_));
 nand2_1 _12116_ (.A(net1239),
    .B(net1699),
    .Y(_07543_));
 or4b_1 _12117_ (.A(net912),
    .B(_07541_),
    .C(_07542_),
    .D_N(_07543_),
    .X(_07544_));
 or3b_1 _12118_ (.A(_07510_),
    .B(_07526_),
    .C_N(_07544_),
    .X(_07545_));
 nand2_1 _12119_ (.A(net1155),
    .B(_07476_),
    .Y(_07546_));
 nor2_1 _12120_ (.A(\digitop_pav2.access_inst.access_ctrl0.ld_key_env_finish_i ),
    .B(_07030_),
    .Y(_07547_));
 nand2_2 _12121_ (.A(_07023_),
    .B(net1063),
    .Y(_07548_));
 or3b_2 _12122_ (.A(net1240),
    .B(_07548_),
    .C_N(_07546_),
    .X(_07549_));
 or2_2 _12123_ (.A(net1240),
    .B(net1017),
    .X(_07550_));
 o21ai_1 _12124_ (.A1(net1154),
    .A2(_07550_),
    .B1(_07549_),
    .Y(_07551_));
 o211a_1 _12125_ (.A1(_07511_),
    .A2(_07551_),
    .B1(_07545_),
    .C1(net963),
    .X(_07552_));
 or3b_1 _12126_ (.A(net1262),
    .B(net201),
    .C_N(\digitop_pav2.access_inst.access_ctrl0.state[10] ),
    .X(_07553_));
 nand2_1 _12127_ (.A(net1260),
    .B(\digitop_pav2.access_inst.access_ctrl0.state[10] ),
    .Y(_07554_));
 and2_1 _12128_ (.A(_07032_),
    .B(\digitop_pav2.access_inst.access_ctrl0.state[11] ),
    .X(_07555_));
 or4_1 _12129_ (.A(\digitop_pav2.access_inst.access_ctrl0.state[2] ),
    .B(\digitop_pav2.access_inst.access_ctrl0.state[14] ),
    .C(\digitop_pav2.access_inst.access_ctrl0.state[18] ),
    .D(_07555_),
    .X(_07556_));
 o21ba_1 _12130_ (.A1(\digitop_pav2.access_inst.access_ctrl0.replay_ok ),
    .A2(_07554_),
    .B1_N(_07556_),
    .X(_07557_));
 a21oi_1 _12131_ (.A1(_07553_),
    .A2(_07557_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.prev_busy ),
    .Y(_07558_));
 a41o_1 _12132_ (.A1(_07021_),
    .A2(\digitop_pav2.access_inst.access_ctrl0.tx_proc_rd_stb_i ),
    .A3(net1037),
    .A4(\digitop_pav2.access_inst.access_ctrl0.state[25] ),
    .B1(_07558_),
    .X(_07559_));
 a21oi_1 _12133_ (.A1(_07026_),
    .A2(net182),
    .B1(_07025_),
    .Y(_07560_));
 nand2_1 _12134_ (.A(net1069),
    .B(_07479_),
    .Y(_07561_));
 and2_1 _12135_ (.A(_07475_),
    .B(net182),
    .X(_07562_));
 o31a_1 _12136_ (.A1(_07560_),
    .A2(_07561_),
    .A3(_07562_),
    .B1(_07491_),
    .X(_07563_));
 nand2_1 _12137_ (.A(\digitop_pav2.access_inst.access_ctrl0.ld_key_env_finish_i ),
    .B(net1063),
    .Y(_07564_));
 nor2_1 _12138_ (.A(net1067),
    .B(_07564_),
    .Y(_07565_));
 or2_1 _12139_ (.A(net1067),
    .B(_07564_),
    .X(_07566_));
 nand2_1 _12140_ (.A(net1148),
    .B(_07475_),
    .Y(_07567_));
 and2_2 _12141_ (.A(\digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt ),
    .B(\digitop_pav2.access_inst.access_ctrl0.ld_dt_stb ),
    .X(_07568_));
 nand2_1 _12142_ (.A(\digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt ),
    .B(\digitop_pav2.access_inst.access_ctrl0.ld_dt_stb ),
    .Y(_07569_));
 or3_1 _12143_ (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[1] ),
    .B(net1049),
    .C(_07569_),
    .X(_07570_));
 a32o_1 _12144_ (.A1(_07479_),
    .A2(_07547_),
    .A3(_07570_),
    .B1(_07567_),
    .B2(_07565_),
    .X(_07571_));
 a21oi_1 _12145_ (.A1(_07026_),
    .A2(_07568_),
    .B1(_07548_),
    .Y(_07572_));
 a21oi_1 _12146_ (.A1(_07026_),
    .A2(net1148),
    .B1(_07547_),
    .Y(_07573_));
 o21ai_1 _12147_ (.A1(_07572_),
    .A2(_07573_),
    .B1(\digitop_pav2.access_inst.access_proc0.proc_crc_check[1] ),
    .Y(_07574_));
 and2_2 _12148_ (.A(net1047),
    .B(\digitop_pav2.access_inst.access_check0.proc_finish1_i ),
    .X(_07575_));
 inv_2 _12149_ (.A(_07575_),
    .Y(_07576_));
 and2b_1 _12150_ (.A_N(\digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt ),
    .B(\digitop_pav2.access_inst.access_ctrl0.ld_dt_stb ),
    .X(_07577_));
 nand2b_1 _12151_ (.A_N(\digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt ),
    .B(\digitop_pav2.access_inst.access_ctrl0.ld_dt_stb ),
    .Y(_07578_));
 nand2_1 _12152_ (.A(_07026_),
    .B(net1033),
    .Y(_07579_));
 nand2_1 _12153_ (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[1] ),
    .B(_07579_),
    .Y(_07580_));
 nand2_1 _12154_ (.A(_07475_),
    .B(net1033),
    .Y(_07581_));
 and3_1 _12155_ (.A(_07493_),
    .B(_07580_),
    .C(_07581_),
    .X(_07582_));
 a221o_1 _12156_ (.A1(_07571_),
    .A2(_07574_),
    .B1(_07582_),
    .B2(_07479_),
    .C1(_07576_),
    .X(_07583_));
 nand2_1 _12157_ (.A(_07026_),
    .B(net1145),
    .Y(_07584_));
 nor2_1 _12158_ (.A(net1145),
    .B(net159),
    .Y(_07585_));
 o2bb2a_1 _12159_ (.A1_N(\digitop_pav2.access_inst.access_proc0.proc_crc_check[1] ),
    .A2_N(_07584_),
    .B1(_07585_),
    .B2(_07476_),
    .X(_07586_));
 o21ai_1 _12160_ (.A1(net1046),
    .A2(_07586_),
    .B1(_07583_),
    .Y(_07587_));
 o32a_1 _12161_ (.A1(_07489_),
    .A2(_07563_),
    .A3(_07587_),
    .B1(_07480_),
    .B2(\digitop_pav2.access_inst.access_proc0.proc_crc_check[1] ),
    .X(_01536_));
 nor2_1 _12162_ (.A(_07026_),
    .B(net182),
    .Y(_07588_));
 a21o_1 _12163_ (.A1(_07026_),
    .A2(net182),
    .B1(_07561_),
    .X(_07589_));
 o21a_1 _12164_ (.A1(_07588_),
    .A2(_07589_),
    .B1(_07491_),
    .X(_07590_));
 nand2_1 _12165_ (.A(net1049),
    .B(_07569_),
    .Y(_07591_));
 nand2_1 _12166_ (.A(net1049),
    .B(_07578_),
    .Y(_07592_));
 a32o_1 _12167_ (.A1(_07493_),
    .A2(_07579_),
    .A3(_07592_),
    .B1(_07591_),
    .B2(_07572_),
    .X(_07593_));
 xor2_1 _12168_ (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[0] ),
    .B(net1147),
    .X(_07594_));
 o2bb2a_1 _12169_ (.A1_N(_07479_),
    .A2_N(_07593_),
    .B1(_07594_),
    .B2(_07566_),
    .X(_07595_));
 o22a_1 _12170_ (.A1(_07026_),
    .A2(net1145),
    .B1(\digitop_pav2.access_inst.access_ctrl0.nvm_busy_i ),
    .B2(_07476_),
    .X(_07596_));
 a21oi_1 _12171_ (.A1(_07584_),
    .A2(_07596_),
    .B1(net1046),
    .Y(_07597_));
 a211o_1 _12172_ (.A1(_07575_),
    .A2(_07595_),
    .B1(_07597_),
    .C1(_07489_),
    .X(_07598_));
 o22a_1 _12173_ (.A1(\digitop_pav2.access_inst.access_proc0.proc_crc_check[0] ),
    .A2(_07480_),
    .B1(_07590_),
    .B2(_07598_),
    .X(_01535_));
 o22a_1 _12174_ (.A1(\digitop_pav2.access_inst.access_ctrl0.crc_init_i ),
    .A2(_07480_),
    .B1(_07489_),
    .B2(net1047),
    .X(_01534_));
 or3_1 _12175_ (.A(net1144),
    .B(_07503_),
    .C(_07564_),
    .X(_07599_));
 nand2_1 _12176_ (.A(net1256),
    .B(net1034),
    .Y(_07600_));
 a31o_1 _12177_ (.A1(net1256),
    .A2(net1034),
    .A3(_07599_),
    .B1(net1260),
    .X(_07601_));
 o31a_1 _12178_ (.A1(net1037),
    .A2(net1238),
    .A3(_07504_),
    .B1(_07601_),
    .X(_07602_));
 nor2_1 _12179_ (.A(_07504_),
    .B(_07509_),
    .Y(_07603_));
 nand2_2 _12180_ (.A(_07503_),
    .B(_07508_),
    .Y(_07604_));
 and3_1 _12181_ (.A(net1065),
    .B(net1151),
    .C(net1319),
    .X(_07605_));
 a41o_1 _12182_ (.A1(_07023_),
    .A2(_07030_),
    .A3(net1069),
    .A4(_07605_),
    .B1(net1260),
    .X(_07606_));
 nand3_2 _12183_ (.A(net1144),
    .B(net1319),
    .C(_07524_),
    .Y(_07607_));
 and2b_1 _12184_ (.A_N(_07606_),
    .B(_07607_),
    .X(_07608_));
 nand2_1 _12185_ (.A(net811),
    .B(_07608_),
    .Y(_07609_));
 a21oi_1 _12186_ (.A1(net1318),
    .A2(_07575_),
    .B1(net1066),
    .Y(_07610_));
 a32o_1 _12187_ (.A1(net1065),
    .A2(net1151),
    .A3(net1318),
    .B1(\digitop_pav2.access_inst.access_ctrl0.state[11] ),
    .B2(net1066),
    .X(_07611_));
 o41a_1 _12188_ (.A1(_07600_),
    .A2(_07609_),
    .A3(_07610_),
    .A4(_07611_),
    .B1(_07602_),
    .X(_07612_));
 o21ai_1 _12189_ (.A1(net964),
    .A2(_07612_),
    .B1(net1190),
    .Y(_07613_));
 or3_1 _12190_ (.A(_07483_),
    .B(net964),
    .C(_07494_),
    .X(_07614_));
 and3b_1 _12191_ (.A_N(_07614_),
    .B(net1238),
    .C(net913),
    .X(_07615_));
 a21o_4 _12192_ (.A1(net1069),
    .A2(_07615_),
    .B1(_07613_),
    .X(_07616_));
 and4_1 _12193_ (.A(net1055),
    .B(net1056),
    .C(net1059),
    .D(net1062),
    .X(_07617_));
 nor2_1 _12194_ (.A(_07052_),
    .B(_07513_),
    .Y(_07618_));
 nand2_1 _12195_ (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[6] ),
    .B(_07512_),
    .Y(_07619_));
 and3_1 _12196_ (.A(net1158),
    .B(net182),
    .C(net1031),
    .X(_07620_));
 and3_1 _12197_ (.A(_07512_),
    .B(net182),
    .C(net1031),
    .X(_07621_));
 and2_1 _12198_ (.A(net1159),
    .B(_07621_),
    .X(_07622_));
 nand2_1 _12199_ (.A(net1052),
    .B(_07622_),
    .Y(_07623_));
 and3b_1 _12200_ (.A_N(net1050),
    .B(net1052),
    .C(_07622_),
    .X(_07624_));
 a21o_1 _12201_ (.A1(net1050),
    .A2(_07623_),
    .B1(_07624_),
    .X(_07625_));
 nor2_1 _12202_ (.A(_07503_),
    .B(net962),
    .Y(_07626_));
 or2_1 _12203_ (.A(_07503_),
    .B(net962),
    .X(_07627_));
 a21o_1 _12204_ (.A1(net1236),
    .A2(net962),
    .B1(_07503_),
    .X(_07628_));
 inv_2 _12205_ (.A(_07628_),
    .Y(_07629_));
 mux2_1 _12206_ (.A0(net1050),
    .A1(_07625_),
    .S(net1037),
    .X(_07630_));
 o21a_2 _12207_ (.A1(\digitop_pav2.access_inst.access_ctrl0.tx_proc_rd_stb_i ),
    .A2(_07558_),
    .B1(net1031),
    .X(_07631_));
 and3_1 _12208_ (.A(net1053),
    .B(_07618_),
    .C(_07631_),
    .X(_07632_));
 xor2_1 _12209_ (.A(net1051),
    .B(_07632_),
    .X(_07633_));
 nor2_1 _12210_ (.A(net1038),
    .B(_07091_),
    .Y(_07634_));
 and3_1 _12211_ (.A(net1061),
    .B(net1069),
    .C(net1151),
    .X(_07635_));
 and3_1 _12212_ (.A(net1069),
    .B(net1151),
    .C(net1031),
    .X(_07636_));
 inv_2 _12213_ (.A(_07636_),
    .Y(_07637_));
 and3_1 _12214_ (.A(net1159),
    .B(_07512_),
    .C(_07636_),
    .X(_07638_));
 nand2_1 _12215_ (.A(net1053),
    .B(_07638_),
    .Y(_07639_));
 and4bb_2 _12216_ (.A_N(net1066),
    .B_N(net1144),
    .C(net1319),
    .D(_07524_),
    .X(_07640_));
 inv_2 _12217_ (.A(_07640_),
    .Y(_07641_));
 nor2_1 _12218_ (.A(_07611_),
    .B(_07640_),
    .Y(_07642_));
 or2_1 _12219_ (.A(_07611_),
    .B(_07640_),
    .X(_07643_));
 xnor2_1 _12220_ (.A(net1051),
    .B(_07639_),
    .Y(_07644_));
 nand2_1 _12221_ (.A(net1061),
    .B(net1150),
    .Y(_07645_));
 nand2_2 _12222_ (.A(net1150),
    .B(net1031),
    .Y(_07646_));
 nor2_1 _12223_ (.A(_07513_),
    .B(_07646_),
    .Y(_07647_));
 inv_2 _12224_ (.A(_07647_),
    .Y(_07648_));
 and3_1 _12225_ (.A(net1053),
    .B(net1159),
    .C(_07647_),
    .X(_07649_));
 xor2_1 _12226_ (.A(net1051),
    .B(_07649_),
    .X(_07650_));
 o22a_1 _12227_ (.A1(_07643_),
    .A2(_07644_),
    .B1(_07650_),
    .B2(_07641_),
    .X(_07651_));
 a21o_1 _12228_ (.A1(_07607_),
    .A2(_07651_),
    .B1(_07606_),
    .X(_07652_));
 or3_2 _12229_ (.A(_07024_),
    .B(net1070),
    .C(net1152),
    .X(_07653_));
 nand2_4 _12230_ (.A(net1233),
    .B(net819),
    .Y(_07654_));
 mux2_1 _12231_ (.A0(_07504_),
    .A1(net1051),
    .S(_07654_),
    .X(_07655_));
 a31o_1 _12232_ (.A1(net1038),
    .A2(_07091_),
    .A3(_07655_),
    .B1(_07024_),
    .X(_07656_));
 nand2_1 _12233_ (.A(net1060),
    .B(net1145),
    .Y(_07657_));
 nand2_1 _12234_ (.A(\digitop_pav2.access_inst.access_ctrl0.crc_en_o ),
    .B(net1032),
    .Y(_07658_));
 or2_1 _12235_ (.A(_07513_),
    .B(_07658_),
    .X(_07659_));
 nor2_1 _12236_ (.A(_07619_),
    .B(_07658_),
    .Y(_07660_));
 nand2_1 _12237_ (.A(net1052),
    .B(_07660_),
    .Y(_07661_));
 a21oi_1 _12238_ (.A1(net1050),
    .A2(_07661_),
    .B1(net1048),
    .Y(_07662_));
 o21ai_1 _12239_ (.A1(net1050),
    .A2(_07661_),
    .B1(_07662_),
    .Y(_07663_));
 or3b_1 _12240_ (.A(_07030_),
    .B(_07655_),
    .C_N(\digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt_ok ),
    .X(_07664_));
 and3_1 _12241_ (.A(net1059),
    .B(net1062),
    .C(net1033),
    .X(_07665_));
 and3_1 _12242_ (.A(net1158),
    .B(net1033),
    .C(net1032),
    .X(_07666_));
 and2_1 _12243_ (.A(net1156),
    .B(_07666_),
    .X(_07667_));
 or3b_1 _12244_ (.A(_07027_),
    .B(_07052_),
    .C_N(_07667_),
    .X(_07668_));
 and2_1 _12245_ (.A(net1050),
    .B(_07668_),
    .X(_07669_));
 nor2_1 _12246_ (.A(net1051),
    .B(_07668_),
    .Y(_07670_));
 nand2_1 _12247_ (.A(_07568_),
    .B(net1031),
    .Y(_07671_));
 nor2_1 _12248_ (.A(_07513_),
    .B(_07671_),
    .Y(_07672_));
 nor2_1 _12249_ (.A(_07619_),
    .B(_07671_),
    .Y(_07673_));
 nand2_1 _12250_ (.A(net1052),
    .B(_07673_),
    .Y(_07674_));
 or2_2 _12251_ (.A(_07030_),
    .B(\digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt_ok ),
    .X(_07675_));
 a21oi_1 _12252_ (.A1(net1050),
    .A2(_07674_),
    .B1(_07675_),
    .Y(_07676_));
 o21ai_1 _12253_ (.A1(net1050),
    .A2(_07674_),
    .B1(_07676_),
    .Y(_07677_));
 o311a_1 _12254_ (.A1(net1064),
    .A2(_07669_),
    .A3(_07670_),
    .B1(net1236),
    .C1(_07510_),
    .X(_07678_));
 a31o_1 _12255_ (.A1(_07664_),
    .A2(_07677_),
    .A3(_07678_),
    .B1(net966),
    .X(_07679_));
 a41o_1 _12256_ (.A1(net1236),
    .A2(net913),
    .A3(_07656_),
    .A4(_07663_),
    .B1(_07679_),
    .X(_07680_));
 nor2_1 _12257_ (.A(net1236),
    .B(net912),
    .Y(_07681_));
 nand2_1 _12258_ (.A(net1262),
    .B(net913),
    .Y(_07682_));
 mux2_1 _12259_ (.A0(_07625_),
    .A1(_07633_),
    .S(net201),
    .X(_07683_));
 o211a_1 _12260_ (.A1(net1236),
    .A2(_07683_),
    .B1(_07652_),
    .C1(net811),
    .X(_07684_));
 a221o_1 _12261_ (.A1(_07629_),
    .A2(_07630_),
    .B1(_07681_),
    .B2(_07625_),
    .C1(_07680_),
    .X(_07685_));
 o22a_1 _12262_ (.A1(net963),
    .A2(_07655_),
    .B1(_07684_),
    .B2(_07685_),
    .X(_07686_));
 mux2_1 _12263_ (.A0(_07686_),
    .A1(net1050),
    .S(_07616_),
    .X(_01533_));
 or2_1 _12264_ (.A(net1052),
    .B(_07622_),
    .X(_07687_));
 nand2_1 _12265_ (.A(_07623_),
    .B(_07687_),
    .Y(_07688_));
 or2_1 _12266_ (.A(net1159),
    .B(_07514_),
    .X(_07689_));
 nor2_1 _12267_ (.A(net1054),
    .B(_07689_),
    .Y(_07690_));
 or3_2 _12268_ (.A(net1054),
    .B(_07542_),
    .C(_07689_),
    .X(_07691_));
 mux2_1 _12269_ (.A0(_07509_),
    .A1(net1052),
    .S(_07654_),
    .X(_07692_));
 inv_2 _12270_ (.A(_07692_),
    .Y(_07693_));
 or2_1 _12271_ (.A(net1052),
    .B(_07660_),
    .X(_07694_));
 nand2_1 _12272_ (.A(_07661_),
    .B(_07694_),
    .Y(_07695_));
 o221a_1 _12273_ (.A1(_07653_),
    .A2(_07693_),
    .B1(_07695_),
    .B2(net1048),
    .C1(net1236),
    .X(_07696_));
 a211o_1 _12274_ (.A1(net1261),
    .A2(_07688_),
    .B1(_07696_),
    .C1(net912),
    .X(_07697_));
 mux2_1 _12275_ (.A0(_07027_),
    .A1(_07688_),
    .S(net1037),
    .X(_07698_));
 o2bb2a_1 _12276_ (.A1_N(net1063),
    .A2_N(net1144),
    .B1(_07673_),
    .B2(net1052),
    .X(_07699_));
 a221o_1 _12277_ (.A1(\digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt_ok ),
    .A2(_07692_),
    .B1(_07699_),
    .B2(_07674_),
    .C1(_07030_),
    .X(_07700_));
 a31o_1 _12278_ (.A1(net1033),
    .A2(net1032),
    .A3(_07618_),
    .B1(net1053),
    .X(_07701_));
 a21oi_1 _12279_ (.A1(_07668_),
    .A2(_07701_),
    .B1(net1064),
    .Y(_07702_));
 or4b_1 _12280_ (.A(net1261),
    .B(_07702_),
    .C(_07511_),
    .D_N(_07700_),
    .X(_07703_));
 or2_1 _12281_ (.A(net1053),
    .B(_07638_),
    .X(_07704_));
 nand2_1 _12282_ (.A(_07639_),
    .B(_07704_),
    .Y(_07705_));
 o21a_1 _12283_ (.A1(_07619_),
    .A2(_07646_),
    .B1(_07027_),
    .X(_07706_));
 o32a_1 _12284_ (.A1(_07641_),
    .A2(_07649_),
    .A3(_07706_),
    .B1(_07705_),
    .B2(_07643_),
    .X(_07707_));
 o211a_1 _12285_ (.A1(_07609_),
    .A2(_07707_),
    .B1(_07703_),
    .C1(net963),
    .X(_07708_));
 o21ai_1 _12286_ (.A1(_07628_),
    .A2(_07698_),
    .B1(_07708_),
    .Y(_07709_));
 or2_1 _12287_ (.A(net1237),
    .B(_07604_),
    .X(_07710_));
 a21oi_1 _12288_ (.A1(_07618_),
    .A2(_07631_),
    .B1(net1053),
    .Y(_07711_));
 or2_1 _12289_ (.A(_07632_),
    .B(_07711_),
    .X(_07712_));
 mux2_1 _12290_ (.A0(_07688_),
    .A1(_07712_),
    .S(net201),
    .X(_07713_));
 o21ai_1 _12291_ (.A1(_07710_),
    .A2(_07713_),
    .B1(_07697_),
    .Y(_07714_));
 o22a_1 _12292_ (.A1(net963),
    .A2(_07692_),
    .B1(_07709_),
    .B2(_07714_),
    .X(_07715_));
 mux2_1 _12293_ (.A0(_07715_),
    .A1(net1052),
    .S(_07616_),
    .X(_01532_));
 a21o_1 _12294_ (.A1(\digitop_pav2.access_inst.access_ctrl0.tx_proc_rd_stb_i ),
    .A2(net201),
    .B1(net182),
    .X(_07716_));
 and3_1 _12295_ (.A(net1058),
    .B(net1062),
    .C(_07716_),
    .X(_07717_));
 and2_1 _12296_ (.A(net1057),
    .B(_07717_),
    .X(_07718_));
 and3_1 _12297_ (.A(net1059),
    .B(net1062),
    .C(_07568_),
    .X(_07719_));
 a21o_1 _12298_ (.A1(net1056),
    .A2(_07719_),
    .B1(net1055),
    .X(_07720_));
 a21o_1 _12299_ (.A1(_07671_),
    .A2(_07720_),
    .B1(_07675_),
    .X(_07721_));
 a21oi_1 _12300_ (.A1(net1056),
    .A2(_07665_),
    .B1(net1055),
    .Y(_07722_));
 a21oi_1 _12301_ (.A1(net1033),
    .A2(net1032),
    .B1(_07722_),
    .Y(_07723_));
 o21a_1 _12302_ (.A1(net1064),
    .A2(_07723_),
    .B1(_07721_),
    .X(_07724_));
 or3_1 _12303_ (.A(net1261),
    .B(_07509_),
    .C(_07724_),
    .X(_07725_));
 o211a_1 _12304_ (.A1(net1054),
    .A2(_07039_),
    .B1(_07504_),
    .C1(_07725_),
    .X(_07726_));
 a21oi_1 _12305_ (.A1(_07681_),
    .A2(_07691_),
    .B1(_07726_),
    .Y(_07727_));
 and3_1 _12306_ (.A(net1058),
    .B(net1060),
    .C(net182),
    .X(_07728_));
 o211ai_1 _12307_ (.A1(_07727_),
    .A2(_07728_),
    .B1(net1032),
    .C1(_07716_),
    .Y(_07729_));
 nor2_1 _12308_ (.A(net1054),
    .B(_07728_),
    .Y(_07730_));
 o21ai_1 _12309_ (.A1(_07727_),
    .A2(_07730_),
    .B1(_07710_),
    .Y(_07731_));
 o211a_1 _12310_ (.A1(net1054),
    .A2(_07718_),
    .B1(_07729_),
    .C1(_07731_),
    .X(_07732_));
 nor2_1 _12311_ (.A(net913),
    .B(_07654_),
    .Y(_07733_));
 mux2_1 _12312_ (.A0(net1054),
    .A1(net1076),
    .S(_07733_),
    .X(_07734_));
 nor2_1 _12313_ (.A(_07029_),
    .B(_07657_),
    .Y(_07735_));
 a21o_1 _12314_ (.A1(net1057),
    .A2(_07735_),
    .B1(net1055),
    .X(_07736_));
 a21o_1 _12315_ (.A1(_07658_),
    .A2(_07736_),
    .B1(net1048),
    .X(_07737_));
 nand2_2 _12316_ (.A(net913),
    .B(_07653_),
    .Y(_07738_));
 nor2_1 _12317_ (.A(net1262),
    .B(_07738_),
    .Y(_07739_));
 o211a_1 _12318_ (.A1(_07024_),
    .A2(_07734_),
    .B1(_07737_),
    .C1(_07739_),
    .X(_07740_));
 and3_1 _12319_ (.A(net1056),
    .B(net1059),
    .C(_07635_),
    .X(_07741_));
 o211a_1 _12320_ (.A1(net1054),
    .A2(_07741_),
    .B1(_07642_),
    .C1(_07637_),
    .X(_07742_));
 nor2_1 _12321_ (.A(_07029_),
    .B(_07645_),
    .Y(_07743_));
 a21o_1 _12322_ (.A1(net1056),
    .A2(_07743_),
    .B1(net1054),
    .X(_07744_));
 a31o_1 _12323_ (.A1(_07640_),
    .A2(_07646_),
    .A3(_07744_),
    .B1(_07742_),
    .X(_07745_));
 a31o_1 _12324_ (.A1(net1236),
    .A2(_07510_),
    .A3(_07724_),
    .B1(net965),
    .X(_07746_));
 a31o_1 _12325_ (.A1(net811),
    .A2(_07608_),
    .A3(_07745_),
    .B1(_07746_),
    .X(_07747_));
 a21o_1 _12326_ (.A1(net1071),
    .A2(_07726_),
    .B1(_07747_),
    .X(_07748_));
 o32a_1 _12327_ (.A1(_07732_),
    .A2(_07740_),
    .A3(_07748_),
    .B1(_07734_),
    .B2(net963),
    .X(_07749_));
 mux2_1 _12328_ (.A0(_07749_),
    .A1(net1054),
    .S(_07616_),
    .X(_01531_));
 xnor2_1 _12329_ (.A(_07028_),
    .B(_07728_),
    .Y(_07750_));
 nor2_1 _12330_ (.A(net1071),
    .B(_07750_),
    .Y(_07751_));
 xnor2_1 _12331_ (.A(_07028_),
    .B(_07719_),
    .Y(_07752_));
 xnor2_1 _12332_ (.A(_07028_),
    .B(_07665_),
    .Y(_07753_));
 o221ai_2 _12333_ (.A1(_07675_),
    .A2(_07752_),
    .B1(_07753_),
    .B2(net1064),
    .C1(_07510_),
    .Y(_07754_));
 a221o_1 _12334_ (.A1(_07028_),
    .A2(net1071),
    .B1(_07628_),
    .B2(_07754_),
    .C1(_07751_),
    .X(_07755_));
 a21oi_1 _12335_ (.A1(net1059),
    .A2(_07635_),
    .B1(net1056),
    .Y(_07756_));
 o21a_1 _12336_ (.A1(_07741_),
    .A2(_07756_),
    .B1(_07642_),
    .X(_07757_));
 xnor2_1 _12337_ (.A(net1056),
    .B(_07743_),
    .Y(_07758_));
 a211o_1 _12338_ (.A1(_07640_),
    .A2(_07758_),
    .B1(_07757_),
    .C1(_07609_),
    .X(_07759_));
 o2111a_1 _12339_ (.A1(net1262),
    .A2(_07754_),
    .B1(_07755_),
    .C1(_07759_),
    .D1(_07488_),
    .X(_07760_));
 a21oi_1 _12340_ (.A1(net1258),
    .A2(net913),
    .B1(_07654_),
    .Y(_07761_));
 a22oi_2 _12341_ (.A1(net1056),
    .A2(_07654_),
    .B1(_07761_),
    .B2(net1078),
    .Y(_07762_));
 xnor2_1 _12342_ (.A(_07028_),
    .B(_07735_),
    .Y(_07763_));
 nor2_1 _12343_ (.A(net1048),
    .B(_07763_),
    .Y(_07764_));
 a211o_1 _12344_ (.A1(net1048),
    .A2(_07762_),
    .B1(_07764_),
    .C1(_07738_),
    .X(_07765_));
 a2bb2o_1 _12345_ (.A1_N(net1237),
    .A2_N(_07750_),
    .B1(_07765_),
    .B2(_07682_),
    .X(_07766_));
 nor2_1 _12346_ (.A(net1057),
    .B(_07717_),
    .Y(_07767_));
 o311a_1 _12347_ (.A1(_07710_),
    .A2(_07718_),
    .A3(_07767_),
    .B1(_07766_),
    .C1(_07760_),
    .X(_07768_));
 a21oi_1 _12348_ (.A1(net965),
    .A2(_07762_),
    .B1(_07768_),
    .Y(_07769_));
 mux2_1 _12349_ (.A0(_07769_),
    .A1(net1057),
    .S(_07616_),
    .X(_01530_));
 nand2_1 _12350_ (.A(net1058),
    .B(_07616_),
    .Y(_07770_));
 a22oi_1 _12351_ (.A1(net1058),
    .A2(_07654_),
    .B1(_07761_),
    .B2(net1080),
    .Y(_07771_));
 and2_1 _12352_ (.A(_07029_),
    .B(_07657_),
    .X(_07772_));
 o21a_1 _12353_ (.A1(_07735_),
    .A2(_07772_),
    .B1(_07024_),
    .X(_07773_));
 a211o_1 _12354_ (.A1(net1048),
    .A2(_07771_),
    .B1(_07773_),
    .C1(_07738_),
    .X(_07774_));
 a21oi_1 _12355_ (.A1(net1060),
    .A2(net182),
    .B1(net1058),
    .Y(_07775_));
 nor2_1 _12356_ (.A(_07728_),
    .B(_07775_),
    .Y(_07776_));
 a21o_1 _12357_ (.A1(net1060),
    .A2(net201),
    .B1(net1058),
    .X(_07777_));
 mux2_1 _12358_ (.A0(_07777_),
    .A1(_07776_),
    .S(_07691_),
    .X(_07778_));
 a2bb2o_1 _12359_ (.A1_N(net1237),
    .A2_N(_07778_),
    .B1(_07774_),
    .B2(_07682_),
    .X(_07779_));
 a21oi_1 _12360_ (.A1(net1062),
    .A2(_07716_),
    .B1(net1058),
    .Y(_07780_));
 xnor2_1 _12361_ (.A(_07029_),
    .B(_07635_),
    .Y(_07781_));
 and2_1 _12362_ (.A(_07029_),
    .B(_07645_),
    .X(_07782_));
 o21ai_1 _12363_ (.A1(_07743_),
    .A2(_07782_),
    .B1(_07640_),
    .Y(_07783_));
 o211a_1 _12364_ (.A1(_07643_),
    .A2(_07781_),
    .B1(_07783_),
    .C1(_07607_),
    .X(_07784_));
 o21ai_1 _12365_ (.A1(_07606_),
    .A2(_07784_),
    .B1(net811),
    .Y(_07785_));
 nor2_1 _12366_ (.A(net1071),
    .B(_07776_),
    .Y(_07786_));
 a21oi_1 _12367_ (.A1(net1062),
    .A2(_07568_),
    .B1(net1059),
    .Y(_07787_));
 or3_1 _12368_ (.A(_07675_),
    .B(_07719_),
    .C(_07787_),
    .X(_07788_));
 a21oi_1 _12369_ (.A1(net1062),
    .A2(net1033),
    .B1(net1059),
    .Y(_07789_));
 or3_1 _12370_ (.A(net1064),
    .B(_07665_),
    .C(_07789_),
    .X(_07790_));
 a31o_1 _12371_ (.A1(net1237),
    .A2(_07788_),
    .A3(_07790_),
    .B1(_07511_),
    .X(_07791_));
 a221o_1 _12372_ (.A1(_07029_),
    .A2(net1071),
    .B1(_07627_),
    .B2(_07791_),
    .C1(_07786_),
    .X(_07792_));
 a21o_1 _12373_ (.A1(_07785_),
    .A2(_07791_),
    .B1(net1261),
    .X(_07793_));
 o311a_1 _12374_ (.A1(_07717_),
    .A2(_07780_),
    .A3(_07785_),
    .B1(_07793_),
    .C1(_07488_),
    .X(_07794_));
 a32o_1 _12375_ (.A1(_07779_),
    .A2(_07792_),
    .A3(_07794_),
    .B1(_07771_),
    .B2(net965),
    .X(_07795_));
 o21ai_1 _12376_ (.A1(_07616_),
    .A2(_07795_),
    .B1(_07770_),
    .Y(_01529_));
 nand2_1 _12377_ (.A(net1061),
    .B(_07616_),
    .Y(_07796_));
 o21a_1 _12378_ (.A1(net1258),
    .A2(_07535_),
    .B1(_07527_),
    .X(_07797_));
 o211a_1 _12379_ (.A1(net1082),
    .A2(_07797_),
    .B1(net818),
    .C1(net1234),
    .X(_07798_));
 a21oi_1 _12380_ (.A1(net1060),
    .A2(_07654_),
    .B1(_07798_),
    .Y(_07799_));
 or2_1 _12381_ (.A(net1060),
    .B(\digitop_pav2.access_inst.access_ctrl0.crc_en_o ),
    .X(_07800_));
 a21oi_1 _12382_ (.A1(_07657_),
    .A2(_07800_),
    .B1(net1048),
    .Y(_07801_));
 a211o_1 _12383_ (.A1(net1048),
    .A2(_07799_),
    .B1(_07801_),
    .C1(_07738_),
    .X(_07802_));
 xor2_1 _12384_ (.A(net1060),
    .B(net182),
    .X(_07803_));
 inv_2 _12385_ (.A(_07803_),
    .Y(_07804_));
 mux2_1 _12386_ (.A0(net202),
    .A1(_07804_),
    .S(_07691_),
    .X(_07805_));
 a22o_1 _12387_ (.A1(_07682_),
    .A2(_07802_),
    .B1(_07805_),
    .B2(net1262),
    .X(_07806_));
 nor2_1 _12388_ (.A(net1061),
    .B(_07634_),
    .Y(_07807_));
 o21ai_1 _12389_ (.A1(_07635_),
    .A2(_07807_),
    .B1(_07642_),
    .Y(_07808_));
 or2_1 _12390_ (.A(net1061),
    .B(net1150),
    .X(_07809_));
 a21o_1 _12391_ (.A1(_07645_),
    .A2(_07809_),
    .B1(_07641_),
    .X(_07810_));
 a31o_1 _12392_ (.A1(_07607_),
    .A2(_07808_),
    .A3(_07810_),
    .B1(_07606_),
    .X(_07811_));
 nand2_1 _12393_ (.A(net811),
    .B(_07811_),
    .Y(_07812_));
 a21oi_1 _12394_ (.A1(net1061),
    .A2(_07716_),
    .B1(_07812_),
    .Y(_07813_));
 o21ai_1 _12395_ (.A1(net1060),
    .A2(_07716_),
    .B1(_07813_),
    .Y(_07814_));
 xnor2_1 _12396_ (.A(net1060),
    .B(_07568_),
    .Y(_07815_));
 nand2b_1 _12397_ (.A_N(net1063),
    .B(\digitop_pav2.access_inst.access_ctrl0.ld_dt_stb ),
    .Y(_07816_));
 a21bo_1 _12398_ (.A1(net1063),
    .A2(net1144),
    .B1_N(_07816_),
    .X(_07817_));
 mux2_1 _12399_ (.A0(_07816_),
    .A1(_07817_),
    .S(_07815_),
    .X(_07818_));
 o21ai_1 _12400_ (.A1(net1262),
    .A2(_07818_),
    .B1(_07510_),
    .Y(_07819_));
 nor2_1 _12401_ (.A(net1061),
    .B(net1037),
    .Y(_07820_));
 a221o_1 _12402_ (.A1(net1037),
    .A2(_07804_),
    .B1(_07819_),
    .B2(_07627_),
    .C1(_07820_),
    .X(_07821_));
 a21o_1 _12403_ (.A1(_07812_),
    .A2(_07819_),
    .B1(net1261),
    .X(_07822_));
 and3_1 _12404_ (.A(net963),
    .B(_07821_),
    .C(_07822_),
    .X(_07823_));
 a32o_1 _12405_ (.A1(_07806_),
    .A2(_07814_),
    .A3(_07823_),
    .B1(_07799_),
    .B2(net964),
    .X(_07824_));
 o21ai_1 _12406_ (.A1(_07616_),
    .A2(_07824_),
    .B1(_07796_),
    .Y(_01528_));
 a31o_1 _12407_ (.A1(net1046),
    .A2(_07490_),
    .A3(_07493_),
    .B1(net1063),
    .X(_01527_));
 a31o_1 _12408_ (.A1(net1046),
    .A2(net1069),
    .A3(_07490_),
    .B1(net1065),
    .X(_01526_));
 o21ai_1 _12409_ (.A1(_07540_),
    .A2(_07559_),
    .B1(net1192),
    .Y(_07825_));
 a22o_1 _12410_ (.A1(net1192),
    .A2(net201),
    .B1(_07825_),
    .B2(\digitop_pav2.access_inst.access_proc0.ctrl_rd_bus ),
    .X(_01525_));
 nor2_1 _12411_ (.A(net1326),
    .B(net1325),
    .Y(_07826_));
 or2_1 _12412_ (.A(net1326),
    .B(net1325),
    .X(_07827_));
 nand2_1 _12413_ (.A(\digitop_pav2.boot_inst.boot_ctrl0.act_state_i ),
    .B(net1322),
    .Y(_07828_));
 mux2_1 _12414_ (.A0(net1771),
    .A1(\digitop_pav2.boot_inst.boot_ctrl0.proc_crc_end_i ),
    .S(_07828_),
    .X(_07829_));
 or4_1 _12415_ (.A(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_crc_en ),
    .B(\digitop_pav2.boot_inst.boot_ctrl0.state[0] ),
    .C(\digitop_pav2.boot_inst.boot_ctrl0.state[2] ),
    .D(net1400),
    .X(_07830_));
 inv_2 _12416_ (.A(_07830_),
    .Y(_07831_));
 or2_2 _12417_ (.A(_07829_),
    .B(_07830_),
    .X(_07832_));
 inv_2 _12418_ (.A(_07832_),
    .Y(_07833_));
 or2_2 _12419_ (.A(_07827_),
    .B(_07832_),
    .X(_07834_));
 nor2_1 _12420_ (.A(_07061_),
    .B(net1317),
    .Y(_07835_));
 nand2_1 _12421_ (.A(\digitop_pav2.boot_inst.boot_ctrl0.proc_boot_end_i ),
    .B(_07828_),
    .Y(_07836_));
 o21ai_2 _12422_ (.A1(\digitop_pav2.boot_inst.boot_ctrl0.act_state_i ),
    .A2(_07835_),
    .B1(net1322),
    .Y(_07837_));
 and2_1 _12423_ (.A(net1771),
    .B(_07837_),
    .X(_07838_));
 or3b_1 _12424_ (.A(_07058_),
    .B(net1783),
    .C_N(_07828_),
    .X(_07839_));
 or4_1 _12425_ (.A(net1755),
    .B(\digitop_pav2.boot_inst.boot_ctrl0.state[0] ),
    .C(\digitop_pav2.boot_inst.boot_ctrl0.state[2] ),
    .D(net1777),
    .X(_07840_));
 and3b_2 _12426_ (.A_N(net1778),
    .B(_07839_),
    .C(_07829_),
    .X(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_replay_o ));
 or2_1 _12427_ (.A(net1400),
    .B(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_replay_o ),
    .X(_07841_));
 or2_2 _12428_ (.A(net1772),
    .B(_07841_),
    .X(_07842_));
 and2b_1 _12429_ (.A_N(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[2] ),
    .B(net1310),
    .X(_07843_));
 or3b_1 _12430_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[1] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[2] ),
    .C_N(net1310),
    .X(_07844_));
 nor2_1 _12431_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[0] ),
    .B(_07844_),
    .Y(_07845_));
 and3b_1 _12432_ (.A_N(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[3] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[2] ),
    .C(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[1] ),
    .X(_07846_));
 nand3b_1 _12433_ (.A_N(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[3] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[2] ),
    .C(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[1] ),
    .Y(_07847_));
 and3_1 _12434_ (.A(_07056_),
    .B(net159),
    .C(_07846_),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_wr_stb ));
 nand2_1 _12435_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[1] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[0] ),
    .Y(_07848_));
 nor2_1 _12436_ (.A(_07056_),
    .B(_07847_),
    .Y(_07849_));
 o31a_1 _12437_ (.A1(_07845_),
    .A2(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_wr_stb ),
    .A3(_07849_),
    .B1(net1482),
    .X(_07850_));
 nand2_2 _12438_ (.A(net1617),
    .B(net1622),
    .Y(_07851_));
 inv_2 _12439_ (.A(net1618),
    .Y(\digitop_pav2.g_auth_obu ));
 and3_2 _12440_ (.A(net715),
    .B(net1626),
    .C(net1629),
    .X(_07852_));
 or3_1 _12441_ (.A(net1050),
    .B(_07497_),
    .C(_07852_),
    .X(_07853_));
 or3b_2 _12442_ (.A(_07853_),
    .B(_07850_),
    .C_N(_07842_),
    .X(_07854_));
 and2b_1 _12443_ (.A_N(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_replay_o ),
    .B(net1772),
    .X(_07855_));
 nand2_2 _12444_ (.A(net1433),
    .B(_07855_),
    .Y(_07856_));
 and2_1 _12445_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[2] ),
    .B(net1269),
    .X(_07857_));
 and2_2 _12446_ (.A(net1269),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[1] ),
    .X(_07858_));
 nand2_1 _12447_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[2] ),
    .B(_07858_),
    .Y(_07859_));
 and2_2 _12448_ (.A(net1268),
    .B(net1178),
    .X(_07860_));
 nand2_1 _12449_ (.A(net1268),
    .B(net1178),
    .Y(_07861_));
 nor2_1 _12450_ (.A(\digitop_pav2.ack_inst.nvm_ack_rd_stb_o ),
    .B(\digitop_pav2.ack_inst.state_ff[1] ),
    .Y(_07862_));
 or2_1 _12451_ (.A(\digitop_pav2.ack_inst.nvm_ack_rd_stb_o ),
    .B(\digitop_pav2.ack_inst.state_ff[1] ),
    .X(_07863_));
 nand2_1 _12452_ (.A(\digitop_pav2.ack_inst.rcnt_ff[0] ),
    .B(\digitop_pav2.ack_inst.rcnt_ff[1] ),
    .Y(_07864_));
 a22o_1 _12453_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[12] ),
    .A2(_07861_),
    .B1(_07863_),
    .B2(_07864_),
    .X(_07865_));
 a2111o_1 _12454_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[6] ),
    .A2(_07859_),
    .B1(_07865_),
    .C1(\digitop_pav2.invent_inst.invent_sel_pav2.state[5] ),
    .D1(_07852_),
    .X(_07866_));
 nor2_1 _12455_ (.A(_07857_),
    .B(_07858_),
    .Y(_07867_));
 or2_1 _12456_ (.A(_07857_),
    .B(_07858_),
    .X(_07868_));
 nand2_1 _12457_ (.A(net1178),
    .B(_07868_),
    .Y(_07869_));
 a22o_1 _12458_ (.A1(net1052),
    .A2(_07498_),
    .B1(_07869_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.state[4] ),
    .X(_07870_));
 or3b_1 _12459_ (.A(_07866_),
    .B(_07870_),
    .C_N(_07856_),
    .X(_07871_));
 and3_1 _12460_ (.A(\digitop_pav2.sec_inst.ld_mem.wctr[2] ),
    .B(\digitop_pav2.sec_inst.ld_mem.round_i ),
    .C(_07852_),
    .X(_07872_));
 a22o_1 _12461_ (.A1(_07498_),
    .A2(_07689_),
    .B1(_07872_),
    .B2(\digitop_pav2.sec_inst.ld_mem.wctr[3] ),
    .X(_07873_));
 and4b_1 _12462_ (.A_N(_07689_),
    .B(_07029_),
    .C(_07028_),
    .D(_07027_),
    .X(_07874_));
 and3_1 _12463_ (.A(net1051),
    .B(net1054),
    .C(_07874_),
    .X(_07875_));
 inv_2 _12464_ (.A(_07875_),
    .Y(_07876_));
 nor2_1 _12465_ (.A(net1618),
    .B(_07872_),
    .Y(_07877_));
 mux2_1 _12466_ (.A0(_07872_),
    .A1(_07877_),
    .S(\digitop_pav2.sec_inst.ld_mem.wctr[3] ),
    .X(_07878_));
 a31o_2 _12467_ (.A1(net1055),
    .A2(_07498_),
    .A3(_07876_),
    .B1(_07878_),
    .X(_07879_));
 or2_2 _12468_ (.A(_07871_),
    .B(_07873_),
    .X(_07880_));
 nor2_1 _12469_ (.A(_07879_),
    .B(_07880_),
    .Y(_07881_));
 or2_1 _12470_ (.A(_07879_),
    .B(_07880_),
    .X(_07882_));
 nor3b_2 _12471_ (.A(_07873_),
    .B(_07879_),
    .C_N(_07871_),
    .Y(_07883_));
 inv_2 _12472_ (.A(_07883_),
    .Y(_07884_));
 nor2_1 _12473_ (.A(net1755),
    .B(_07058_),
    .Y(_07885_));
 a211oi_1 _12474_ (.A1(_07838_),
    .A2(net1756),
    .B1(_07841_),
    .C1(_07827_),
    .Y(_07886_));
 nor2_1 _12475_ (.A(_07850_),
    .B(_07875_),
    .Y(_07887_));
 or2_1 _12476_ (.A(\digitop_pav2.ack_inst.rcnt_ff[0] ),
    .B(_07062_),
    .X(_07888_));
 nor2_1 _12477_ (.A(_07862_),
    .B(_07888_),
    .Y(_07889_));
 or3_1 _12478_ (.A(net1057),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.state[5] ),
    .C(_07889_),
    .X(_07890_));
 and3_1 _12479_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[6] ),
    .B(_07859_),
    .C(_07868_),
    .X(_07891_));
 nor2_1 _12480_ (.A(net1178),
    .B(_07859_),
    .Y(_07892_));
 a21o_1 _12481_ (.A1(\digitop_pav2.sec_inst.en_ld_data ),
    .A2(\digitop_pav2.sec_inst.ld_mem.round_i ),
    .B1(\digitop_pav2.sec_inst.ld_mem.wctr[2] ),
    .X(_07893_));
 a221o_1 _12482_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[12] ),
    .A2(_07892_),
    .B1(_07893_),
    .B2(_07877_),
    .C1(_07891_),
    .X(_07894_));
 a311o_1 _12483_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[4] ),
    .A2(_07860_),
    .A3(_07867_),
    .B1(_07890_),
    .C1(_07894_),
    .X(_07895_));
 or4b_2 _12484_ (.A(_07497_),
    .B(_07895_),
    .C(net1757),
    .D_N(_07887_),
    .X(_07896_));
 o21bai_1 _12485_ (.A1(net1761),
    .A2(net1756),
    .B1_N(net1752),
    .Y(_07897_));
 o211ai_4 _12486_ (.A1(\digitop_pav2.boot_inst.boot_ctrl0.act_state_i ),
    .A2(\digitop_pav2.acc_activate ),
    .B1(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_replay_o ),
    .C1(net1322),
    .Y(_07898_));
 inv_2 _12487_ (.A(net1030),
    .Y(_07899_));
 nor2_1 _12488_ (.A(_07860_),
    .B(_07868_),
    .Y(_07900_));
 nand2_1 _12489_ (.A(_07861_),
    .B(_07867_),
    .Y(_07901_));
 nor2_1 _12490_ (.A(_07892_),
    .B(_07900_),
    .Y(_07902_));
 a21o_1 _12491_ (.A1(net1030),
    .A2(_07900_),
    .B1(_07892_),
    .X(_07903_));
 nand2_1 _12492_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[4] ),
    .B(_07903_),
    .Y(_07904_));
 nand2_1 _12493_ (.A(\digitop_pav2.ack_inst.rcnt_ff[0] ),
    .B(_07062_),
    .Y(_07905_));
 a32o_1 _12494_ (.A1(\digitop_pav2.ack_inst.rcnt_ff[0] ),
    .A2(_07062_),
    .A3(_07863_),
    .B1(net1008),
    .B2(\digitop_pav2.sec_inst.ld_mem.wctr[0] ),
    .X(_07906_));
 nand2_1 _12495_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[6] ),
    .B(_07867_),
    .Y(_07907_));
 or4b_1 _12496_ (.A(net1062),
    .B(_07497_),
    .C(_07906_),
    .D_N(_07907_),
    .X(_07908_));
 and3_1 _12497_ (.A(_07859_),
    .B(_07861_),
    .C(_07868_),
    .X(_07909_));
 a21oi_1 _12498_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[12] ),
    .A2(_07909_),
    .B1(_07908_),
    .Y(_07910_));
 o211a_1 _12499_ (.A1(net1761),
    .A2(_07842_),
    .B1(_07887_),
    .C1(_07910_),
    .X(_07911_));
 o211ai_4 _12500_ (.A1(_07856_),
    .A2(_07897_),
    .B1(_07904_),
    .C1(net1762),
    .Y(_07912_));
 a221o_1 _12501_ (.A1(\digitop_pav2.sec_inst.ld_mem.wctr[1] ),
    .A2(net1008),
    .B1(_07863_),
    .B2(_07062_),
    .C1(net1058),
    .X(_07913_));
 or3b_1 _12502_ (.A(net1178),
    .B(_07867_),
    .C_N(\digitop_pav2.invent_inst.invent_sel_pav2.state[4] ),
    .X(_07914_));
 a31o_1 _12503_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[12] ),
    .A2(_07859_),
    .A3(_07861_),
    .B1(_07913_),
    .X(_07915_));
 and3_1 _12504_ (.A(_07498_),
    .B(_07887_),
    .C(_07907_),
    .X(_07916_));
 and3b_1 _12505_ (.A_N(_07915_),
    .B(_07916_),
    .C(_07914_),
    .X(_07917_));
 o221a_1 _12506_ (.A1(net1752),
    .A2(_07842_),
    .B1(_07856_),
    .B2(_07826_),
    .C1(_07917_),
    .X(_07918_));
 o221ai_4 _12507_ (.A1(net1325),
    .A2(net1773),
    .B1(_07856_),
    .B2(_07826_),
    .C1(_07917_),
    .Y(_07919_));
 o21ai_1 _12508_ (.A1(net1763),
    .A2(net1774),
    .B1(_07896_),
    .Y(_07920_));
 a21oi_1 _12509_ (.A1(_07879_),
    .A2(_07920_),
    .B1(_07880_),
    .Y(_07921_));
 o22a_1 _12510_ (.A1(_07854_),
    .A2(_07881_),
    .B1(_07883_),
    .B2(_07921_),
    .X(_07922_));
 or2_1 _12511_ (.A(_07896_),
    .B(_07919_),
    .X(_07923_));
 and4b_1 _12512_ (.A_N(_07854_),
    .B(_07883_),
    .C(_07920_),
    .D(_07923_),
    .X(_07924_));
 nor2_1 _12513_ (.A(_07922_),
    .B(_07924_),
    .Y(_07925_));
 or3_1 _12514_ (.A(_07854_),
    .B(_07884_),
    .C(_07923_),
    .X(_07926_));
 or2_1 _12515_ (.A(net1763),
    .B(_07926_),
    .X(_07927_));
 o21a_1 _12516_ (.A1(net1763),
    .A2(_07925_),
    .B1(_07927_),
    .X(_07928_));
 nand2_1 _12517_ (.A(_07925_),
    .B(_07927_),
    .Y(_07929_));
 and2_1 _12518_ (.A(\digitop_pav2.memctrl_inst.nvm_wr_en_i ),
    .B(_07929_),
    .X(_07930_));
 o21a_2 _12519_ (.A1(\digitop_pav2.memctrl_inst.nvm_rd_en_i ),
    .A2(\digitop_pav2.memctrl_inst.nvm_wr_en_i ),
    .B1(_07929_),
    .X(_07931_));
 and2b_1 _12520_ (.A_N(_07926_),
    .B(net1763),
    .X(_07932_));
 xnor2_1 _12521_ (.A(\digitop_pav2.memctrl_inst.flops_0x081[3] ),
    .B(net1125),
    .Y(_07933_));
 xor2_1 _12522_ (.A(\digitop_pav2.memctrl_inst.flops_0x081[7] ),
    .B(net1111),
    .X(_07934_));
 a2bb2o_1 _12523_ (.A1_N(\digitop_pav2.memctrl_inst.flops_0x081[0] ),
    .A2_N(_07073_),
    .B1(\digitop_pav2.memctrl_inst.flops_0x081[13] ),
    .B2(_07082_),
    .X(_07935_));
 a22o_1 _12524_ (.A1(\digitop_pav2.memctrl_inst.flops_0x081[6] ),
    .A2(_07078_),
    .B1(\digitop_pav2.memctrl_inst.flops_0x081[12] ),
    .B2(net1035),
    .X(_07936_));
 xor2_1 _12525_ (.A(net1084),
    .B(\digitop_pav2.memctrl_inst.flops_0x081[15] ),
    .X(_07937_));
 xor2_1 _12526_ (.A(\digitop_pav2.memctrl_inst.flops_0x081[11] ),
    .B(net1096),
    .X(_07938_));
 xor2_1 _12527_ (.A(\digitop_pav2.memctrl_inst.flops_0x081[9] ),
    .B(net1103),
    .X(_07939_));
 o221ai_1 _12528_ (.A1(\digitop_pav2.memctrl_inst.flops_0x081[12] ),
    .A2(net1035),
    .B1(\digitop_pav2.memctrl_inst.flops_0x081[13] ),
    .B2(_07082_),
    .C1(_07933_),
    .Y(_07940_));
 xor2_1 _12529_ (.A(\digitop_pav2.memctrl_inst.flops_0x081[8] ),
    .B(net1107),
    .X(_07941_));
 xor2_1 _12530_ (.A(\digitop_pav2.memctrl_inst.flops_0x081[10] ),
    .B(net1100),
    .X(_07942_));
 o22a_1 _12531_ (.A1(\digitop_pav2.memctrl_inst.flops_0x081[2] ),
    .A2(_07075_),
    .B1(\digitop_pav2.memctrl_inst.flops_0x081[4] ),
    .B2(_07076_),
    .X(_07943_));
 xnor2_1 _12532_ (.A(\digitop_pav2.memctrl_inst.flops_0x081[1] ),
    .B(net1131),
    .Y(_07944_));
 a221o_1 _12533_ (.A1(\digitop_pav2.memctrl_inst.flops_0x081[0] ),
    .A2(_07073_),
    .B1(\digitop_pav2.memctrl_inst.flops_0x081[14] ),
    .B2(_07083_),
    .C1(_07935_),
    .X(_07945_));
 o221ai_1 _12534_ (.A1(_07074_),
    .A2(net1128),
    .B1(\digitop_pav2.memctrl_inst.flops_0x081[6] ),
    .B2(_07078_),
    .C1(_07943_),
    .Y(_07946_));
 o221ai_1 _12535_ (.A1(\digitop_pav2.memctrl_inst.flops_0x081[5] ),
    .A2(_07077_),
    .B1(\digitop_pav2.memctrl_inst.flops_0x081[14] ),
    .B2(_07083_),
    .C1(_07944_),
    .Y(_07947_));
 a221o_1 _12536_ (.A1(\digitop_pav2.memctrl_inst.flops_0x081[4] ),
    .A2(_07076_),
    .B1(\digitop_pav2.memctrl_inst.flops_0x081[5] ),
    .B2(_07077_),
    .C1(_07936_),
    .X(_07948_));
 or4_1 _12537_ (.A(_07945_),
    .B(_07946_),
    .C(_07947_),
    .D(_07948_),
    .X(_07949_));
 or4_1 _12538_ (.A(_07934_),
    .B(_07938_),
    .C(_07939_),
    .D(_07941_),
    .X(_07950_));
 or4_1 _12539_ (.A(_07937_),
    .B(_07940_),
    .C(_07942_),
    .D(_07950_),
    .X(_07951_));
 nand2_1 _12540_ (.A(\digitop_pav2.memctrl_inst.nvm_wr_en_i ),
    .B(_07932_),
    .Y(_07952_));
 inv_2 _12541_ (.A(net151),
    .Y(_07953_));
 or3_1 _12542_ (.A(_07896_),
    .B(net1763),
    .C(net1753),
    .X(_07954_));
 o211a_1 _12543_ (.A1(_07949_),
    .A2(_07951_),
    .B1(\digitop_pav2.memctrl_inst.nvm_rd_en_i ),
    .C1(_07932_),
    .X(_07955_));
 and4bb_1 _12544_ (.A_N(_07880_),
    .B_N(_07954_),
    .C(_07854_),
    .D(_07879_),
    .X(_07956_));
 a21o_1 _12545_ (.A1(\digitop_pav2.memctrl_inst.nvm_rd_en_i ),
    .A2(_07956_),
    .B1(net149),
    .X(_07957_));
 a211o_1 _12546_ (.A1(\digitop_pav2.memctrl_inst.nvm_wr_en_i ),
    .A2(_07956_),
    .B1(_07957_),
    .C1(_07953_),
    .X(_07958_));
 or3_4 _12547_ (.A(net1634),
    .B(_07931_),
    .C(_07958_),
    .X(\digitop_pav2.access_inst.access_ctrl0.nvm_busy_i ));
 nor2_1 _12548_ (.A(\digitop_pav2.access_inst.access_ctrl0.nvm_busy_i ),
    .B(net1204),
    .Y(_07959_));
 nand2_4 _12549_ (.A(_07237_),
    .B(net1190),
    .Y(_07960_));
 o21a_1 _12550_ (.A1(\digitop_pav2.access_inst.access_ctrl0.prev_busy ),
    .A2(net1191),
    .B1(_07960_),
    .X(_01524_));
 nand2_1 _12551_ (.A(\digitop_pav2.access_inst.access_ctrl0.tx_proc_rd_stb_i ),
    .B(net1192),
    .Y(_07961_));
 mux2_1 _12552_ (.A0(net201),
    .A1(\digitop_pav2.access_inst.access_proc0.ctrl_rd_bus_res ),
    .S(_07961_),
    .X(_01523_));
 o31a_1 _12553_ (.A1(\digitop_pav2.access_inst.access_ctrl0.state[9] ),
    .A2(\digitop_pav2.access_inst.access_ctrl0.state[24] ),
    .A3(\digitop_pav2.access_inst.access_ctrl0.state[23] ),
    .B1(_07031_),
    .X(_07962_));
 or4_1 _12554_ (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[4] ),
    .B(\digitop_pav2.access_inst.access_proc0.proc_crc_check[3] ),
    .C(_07478_),
    .D(_07481_),
    .X(_07963_));
 nor2_1 _12555_ (.A(_07483_),
    .B(_07963_),
    .Y(_07964_));
 a41o_1 _12556_ (.A1(_07495_),
    .A2(_07565_),
    .A3(net1016),
    .A4(_07964_),
    .B1(net1067),
    .X(_01522_));
 nand3_1 _12557_ (.A(net1702),
    .B(\digitop_pav2.access_inst.access_check0.mem_sign_check_i ),
    .C(net1018),
    .Y(_07965_));
 mux2_1 _12558_ (.A0(_07053_),
    .A1(\digitop_pav2.access_inst.access_check0.wcnt_check_zero ),
    .S(_07965_),
    .X(_01521_));
 nor2_1 _12559_ (.A(_07104_),
    .B(net1207),
    .Y(_07966_));
 or2_1 _12560_ (.A(\digitop_pav2.access_inst.access_check0.pc_lock_check_sync_o ),
    .B(_07966_),
    .X(_01520_));
 nand2_1 _12561_ (.A(net1239),
    .B(_07966_),
    .Y(_07967_));
 nand4_1 _12562_ (.A(net1699),
    .B(net1081),
    .C(_07531_),
    .D(_07534_),
    .Y(_07968_));
 or4_1 _12563_ (.A(net1079),
    .B(net912),
    .C(_07967_),
    .D(_07968_),
    .X(_07969_));
 a21bo_1 _12564_ (.A1(\digitop_pav2.access_inst.access_check0.pc_invalid_o ),
    .A2(_07967_),
    .B1_N(_07969_),
    .X(_01519_));
 and2_1 _12565_ (.A(\digitop_pav2.access_inst.access_check0.mem_sign_check_i ),
    .B(net1192),
    .X(_07970_));
 nor2_1 _12566_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[2] ),
    .B(net1077),
    .Y(_07971_));
 xor2_1 _12567_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[3] ),
    .B(net1076),
    .X(_07972_));
 xnor2_1 _12568_ (.A(_07971_),
    .B(_07972_),
    .Y(_07973_));
 or2_1 _12569_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[1] ),
    .B(net1079),
    .X(_07974_));
 and2_1 _12570_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[2] ),
    .B(net1077),
    .X(_07975_));
 o21ai_1 _12571_ (.A1(_07971_),
    .A2(_07975_),
    .B1(_07974_),
    .Y(_07976_));
 or3_1 _12572_ (.A(_07971_),
    .B(_07974_),
    .C(_07975_),
    .X(_07977_));
 nand2_1 _12573_ (.A(_07976_),
    .B(_07977_),
    .Y(_07978_));
 nand2_1 _12574_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[1] ),
    .B(net1079),
    .Y(_07979_));
 nor2_1 _12575_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[0] ),
    .B(net1082),
    .Y(_07980_));
 a21o_1 _12576_ (.A1(_07974_),
    .A2(_07979_),
    .B1(_07980_),
    .X(_07981_));
 or2_1 _12577_ (.A(_07978_),
    .B(_07981_),
    .X(_07982_));
 a21o_1 _12578_ (.A1(_07976_),
    .A2(_07982_),
    .B1(_07973_),
    .X(_07983_));
 and2_1 _12579_ (.A(_07389_),
    .B(_07395_),
    .X(_07984_));
 nand2_1 _12580_ (.A(_07389_),
    .B(_07395_),
    .Y(_07985_));
 a31oi_1 _12581_ (.A1(_07973_),
    .A2(_07976_),
    .A3(_07982_),
    .B1(_07985_),
    .Y(_07986_));
 or2_1 _12582_ (.A(\digitop_pav2.access_inst.access_check0.error_wordcnt_i ),
    .B(\digitop_pav2.access_inst.access_check0.error_word_cnt_ptr ),
    .X(_07987_));
 a221o_1 _12583_ (.A1(net1076),
    .A2(_07985_),
    .B1(_07986_),
    .B2(_07983_),
    .C1(_07987_),
    .X(_07988_));
 nor2_1 _12584_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[5] ),
    .B(net1073),
    .Y(_07989_));
 xor2_1 _12585_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[6] ),
    .B(net1072),
    .X(_07990_));
 or2_1 _12586_ (.A(_07989_),
    .B(_07990_),
    .X(_07991_));
 o21a_1 _12587_ (.A1(_07971_),
    .A2(_07972_),
    .B1(_07983_),
    .X(_07992_));
 nor2_1 _12588_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[4] ),
    .B(net1074),
    .Y(_07993_));
 and2_1 _12589_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[5] ),
    .B(net1073),
    .X(_07994_));
 or2_1 _12590_ (.A(_07989_),
    .B(_07994_),
    .X(_07995_));
 inv_2 _12591_ (.A(_07995_),
    .Y(_07996_));
 xor2_1 _12592_ (.A(_07993_),
    .B(_07995_),
    .X(_07997_));
 and2_1 _12593_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[4] ),
    .B(net1074),
    .X(_07998_));
 o22a_1 _12594_ (.A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[3] ),
    .A2(net1075),
    .B1(_07993_),
    .B2(_07998_),
    .X(_07999_));
 or4_1 _12595_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[3] ),
    .B(net1076),
    .C(_07993_),
    .D(_07998_),
    .X(_08000_));
 or4b_1 _12596_ (.A(_07992_),
    .B(_07997_),
    .C(_07999_),
    .D_N(_08000_),
    .X(_08001_));
 nand2b_1 _12597_ (.A_N(_07997_),
    .B(_07999_),
    .Y(_08002_));
 o211a_1 _12598_ (.A1(_07993_),
    .A2(_07996_),
    .B1(_08001_),
    .C1(_08002_),
    .X(_08003_));
 nand2_1 _12599_ (.A(_07989_),
    .B(_07990_),
    .Y(_08004_));
 and2_1 _12600_ (.A(_07991_),
    .B(_08004_),
    .X(_08005_));
 inv_2 _12601_ (.A(_08005_),
    .Y(_08006_));
 o21ai_1 _12602_ (.A1(_08003_),
    .A2(_08006_),
    .B1(_07991_),
    .Y(_08007_));
 mux2_1 _12603_ (.A0(_07539_),
    .A1(_08007_),
    .S(_07389_),
    .X(_08008_));
 o21a_1 _12604_ (.A1(_07396_),
    .A2(_08008_),
    .B1(net1072),
    .X(_08009_));
 xnor2_1 _12605_ (.A(_08003_),
    .B(_08005_),
    .Y(_08010_));
 a21o_1 _12606_ (.A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[6] ),
    .A2(_08007_),
    .B1(_08010_),
    .X(_08011_));
 o211a_1 _12607_ (.A1(_07389_),
    .A2(_07539_),
    .B1(_08011_),
    .C1(_07395_),
    .X(_08012_));
 o21ai_1 _12608_ (.A1(_07996_),
    .A2(_08000_),
    .B1(_08002_),
    .Y(_08013_));
 nand2_1 _12609_ (.A(_07992_),
    .B(_08013_),
    .Y(_08014_));
 and3_1 _12610_ (.A(_07984_),
    .B(_08001_),
    .C(_08014_),
    .X(_08015_));
 a2111o_1 _12611_ (.A1(_07530_),
    .A2(_07985_),
    .B1(_08009_),
    .C1(_08012_),
    .D1(_08015_),
    .X(_08016_));
 a21o_1 _12612_ (.A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[0] ),
    .A2(_07539_),
    .B1(_07985_),
    .X(_08017_));
 a22o_1 _12613_ (.A1(_07980_),
    .A2(_07984_),
    .B1(_08017_),
    .B2(net1081),
    .X(_08018_));
 nand2_1 _12614_ (.A(_07981_),
    .B(_07984_),
    .Y(_08019_));
 a31oi_1 _12615_ (.A1(_07974_),
    .A2(_07979_),
    .A3(_07980_),
    .B1(_08019_),
    .Y(_08020_));
 a21o_1 _12616_ (.A1(net1080),
    .A2(_07985_),
    .B1(_08020_),
    .X(_08021_));
 and2_1 _12617_ (.A(net1077),
    .B(_07985_),
    .X(_08022_));
 nand2_1 _12618_ (.A(_07978_),
    .B(_07981_),
    .Y(_08023_));
 a31o_1 _12619_ (.A1(_07982_),
    .A2(_07984_),
    .A3(_08023_),
    .B1(_08022_),
    .X(_08024_));
 o21a_1 _12620_ (.A1(_08018_),
    .A2(_08021_),
    .B1(_08024_),
    .X(_08025_));
 o21a_1 _12621_ (.A1(_08016_),
    .A2(_08025_),
    .B1(_07527_),
    .X(_08026_));
 o21a_1 _12622_ (.A1(_07988_),
    .A2(_08026_),
    .B1(_07511_),
    .X(_08027_));
 a211o_1 _12623_ (.A1(_08018_),
    .A2(_08021_),
    .B1(_08024_),
    .C1(_07987_),
    .X(_08028_));
 a21oi_1 _12624_ (.A1(_07988_),
    .A2(_08028_),
    .B1(_08016_),
    .Y(_08029_));
 and4b_1 _12625_ (.A_N(net1075),
    .B(net1077),
    .C(net1079),
    .D(net1081),
    .X(_08030_));
 a21o_1 _12626_ (.A1(net1075),
    .A2(_07535_),
    .B1(_08030_),
    .X(_08031_));
 and2_1 _12627_ (.A(net1077),
    .B(net1075),
    .X(_08032_));
 nand2_1 _12628_ (.A(_07531_),
    .B(_08031_),
    .Y(_08033_));
 and4b_1 _12629_ (.A_N(_07533_),
    .B(_08032_),
    .C(net1694),
    .D(_07531_),
    .X(_08034_));
 nor2_2 _12630_ (.A(_07069_),
    .B(_08033_),
    .Y(_08035_));
 or4_1 _12631_ (.A(_07511_),
    .B(_08029_),
    .C(_08034_),
    .D(_08035_),
    .X(_08036_));
 nand2_1 _12632_ (.A(_07970_),
    .B(_08036_),
    .Y(_08037_));
 o22a_1 _12633_ (.A1(\digitop_pav2.access_inst.access_check0.error_word_cnt_ptr ),
    .A2(_07970_),
    .B1(_08027_),
    .B2(_08037_),
    .X(_01517_));
 nand2_1 _12634_ (.A(\digitop_pav2.access_inst.access_check0.wr_lock_ck_i ),
    .B(net1193),
    .Y(_08038_));
 o21a_1 _12635_ (.A1(net1149),
    .A2(net1151),
    .B1(net1193),
    .X(_08039_));
 and2b_1 _12636_ (.A_N(_08039_),
    .B(_08038_),
    .X(_08040_));
 or2_1 _12637_ (.A(\digitop_pav2.access_inst.access_check0.ctrl_wcknzero_ck ),
    .B(_08040_),
    .X(_08041_));
 nand2_1 _12638_ (.A(net1073),
    .B(net1074),
    .Y(_08042_));
 nand2_1 _12639_ (.A(_07530_),
    .B(_08042_),
    .Y(_08043_));
 mux2_1 _12640_ (.A0(\digitop_pav2.access_inst.access_proc0.ctrl_rd_bus ),
    .A1(\digitop_pav2.access_inst.access_proc0.ctrl_rd_bus_res ),
    .S(_08043_),
    .X(_08044_));
 o211ai_4 _12641_ (.A1(_07509_),
    .A2(_08044_),
    .B1(net963),
    .C1(_07503_),
    .Y(_08045_));
 nand2_1 _12642_ (.A(net1256),
    .B(net1145),
    .Y(_08046_));
 a31o_1 _12643_ (.A1(net1256),
    .A2(\digitop_pav2.access_inst.access_ctrl0.crc_en_o ),
    .A3(net201),
    .B1(\digitop_pav2.access_inst.access_proc0.ctrl_rd_bus ),
    .X(_08047_));
 inv_2 _12644_ (.A(_08047_),
    .Y(_08048_));
 a21o_1 _12645_ (.A1(_07509_),
    .A2(_08048_),
    .B1(_08045_),
    .X(_08049_));
 nand2_2 _12646_ (.A(net1086),
    .B(net180),
    .Y(_08050_));
 inv_2 _12647_ (.A(_08050_),
    .Y(_08051_));
 and2_1 _12648_ (.A(net1120),
    .B(net179),
    .X(_08052_));
 nand2_2 _12649_ (.A(net1118),
    .B(net180),
    .Y(_08053_));
 and2_2 _12650_ (.A(net1114),
    .B(net179),
    .X(_08054_));
 nand2_2 _12651_ (.A(net1114),
    .B(net179),
    .Y(_08055_));
 and2_1 _12652_ (.A(net1132),
    .B(net179),
    .X(_08056_));
 nand2_2 _12653_ (.A(net1132),
    .B(net181),
    .Y(_08057_));
 and2_1 _12654_ (.A(net1130),
    .B(net180),
    .X(_08058_));
 nand2_2 _12655_ (.A(net1127),
    .B(net180),
    .Y(_08059_));
 nand2_2 _12656_ (.A(net1135),
    .B(net180),
    .Y(_08060_));
 and2_1 _12657_ (.A(net1106),
    .B(net179),
    .X(_08061_));
 nand2_2 _12658_ (.A(net1106),
    .B(net180),
    .Y(_08062_));
 o21ai_1 _12659_ (.A1(net1097),
    .A2(_08047_),
    .B1(net913),
    .Y(_08063_));
 o2bb2a_4 _12660_ (.A1_N(net1097),
    .A2_N(_08045_),
    .B1(_08063_),
    .B2(net964),
    .X(_08064_));
 inv_2 _12661_ (.A(_08064_),
    .Y(_08065_));
 o21ai_1 _12662_ (.A1(net1095),
    .A2(_08047_),
    .B1(net913),
    .Y(_08066_));
 o2bb2a_4 _12663_ (.A1_N(net1094),
    .A2_N(_08045_),
    .B1(_08066_),
    .B2(net964),
    .X(_08067_));
 inv_2 _12664_ (.A(_08067_),
    .Y(_08068_));
 and2_1 _12665_ (.A(net1110),
    .B(net179),
    .X(_08069_));
 nand2_2 _12666_ (.A(net1107),
    .B(net180),
    .Y(_08070_));
 xnor2_1 _12667_ (.A(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[8] ),
    .B(_08070_),
    .Y(_08071_));
 nand2_2 _12668_ (.A(net1090),
    .B(net180),
    .Y(_08072_));
 inv_2 _12669_ (.A(_08072_),
    .Y(_08073_));
 and2_1 _12670_ (.A(net1102),
    .B(net179),
    .X(_08074_));
 nand2_2 _12671_ (.A(net1099),
    .B(net180),
    .Y(_08075_));
 xnor2_1 _12672_ (.A(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[10] ),
    .B(_08075_),
    .Y(_08076_));
 and2_1 _12673_ (.A(net1126),
    .B(net181),
    .X(_08077_));
 nand2_2 _12674_ (.A(net1126),
    .B(net181),
    .Y(_08078_));
 xnor2_1 _12675_ (.A(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[3] ),
    .B(_08078_),
    .Y(_08079_));
 and2_1 _12676_ (.A(net1123),
    .B(net179),
    .X(_08080_));
 nand2_2 _12677_ (.A(net1121),
    .B(net181),
    .Y(_08081_));
 and2_1 _12678_ (.A(net1117),
    .B(net179),
    .X(_08082_));
 nand2_2 _12679_ (.A(net1117),
    .B(net181),
    .Y(_08083_));
 nand2_2 _12680_ (.A(net1089),
    .B(net179),
    .Y(_08084_));
 inv_2 _12681_ (.A(_08084_),
    .Y(_08085_));
 xnor2_1 _12682_ (.A(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[14] ),
    .B(_08084_),
    .Y(_08086_));
 a2bb2o_1 _12683_ (.A1_N(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[4] ),
    .A2_N(_08081_),
    .B1(_08059_),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[2] ),
    .X(_08087_));
 a2bb2o_1 _12684_ (.A1_N(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[0] ),
    .A2_N(_08060_),
    .B1(_08055_),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[7] ),
    .X(_08088_));
 a22o_1 _12685_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[1] ),
    .A2(_08057_),
    .B1(_08081_),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[4] ),
    .X(_08089_));
 o22ai_1 _12686_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[7] ),
    .A2(_08055_),
    .B1(_08059_),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[2] ),
    .Y(_08090_));
 a221o_1 _12687_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[15] ),
    .A2(_08050_),
    .B1(_08062_),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[9] ),
    .C1(_08076_),
    .X(_08091_));
 a2bb2o_1 _12688_ (.A1_N(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[1] ),
    .A2_N(_08057_),
    .B1(_08060_),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[0] ),
    .X(_08092_));
 a221o_1 _12689_ (.A1(_07102_),
    .A2(_08061_),
    .B1(_08083_),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[6] ),
    .C1(_08092_),
    .X(_08093_));
 or4_1 _12690_ (.A(_08089_),
    .B(_08090_),
    .C(_08091_),
    .D(_08093_),
    .X(_08094_));
 a2bb2o_1 _12691_ (.A1_N(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[15] ),
    .A2_N(_08050_),
    .B1(_08053_),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[5] ),
    .X(_08095_));
 o22ai_1 _12692_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[5] ),
    .A2(_08053_),
    .B1(_08083_),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[6] ),
    .Y(_08096_));
 a2bb2o_1 _12693_ (.A1_N(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[11] ),
    .A2_N(_08064_),
    .B1(_08072_),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[13] ),
    .X(_08097_));
 xnor2_1 _12694_ (.A(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[12] ),
    .B(_08067_),
    .Y(_08098_));
 a211o_1 _12695_ (.A1(_07103_),
    .A2(_08073_),
    .B1(_08097_),
    .C1(_08098_),
    .X(_08099_));
 a2111o_1 _12696_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[11] ),
    .A2(_08064_),
    .B1(_08079_),
    .C1(_08095_),
    .D1(_08096_),
    .X(_08100_));
 or4_1 _12697_ (.A(_08071_),
    .B(_08086_),
    .C(_08087_),
    .D(_08088_),
    .X(_08101_));
 or4_1 _12698_ (.A(_08094_),
    .B(_08099_),
    .C(_08100_),
    .D(_08101_),
    .X(_08102_));
 xnor2_1 _12699_ (.A(\digitop_pav2.access_inst.access_check0.fg_i[8] ),
    .B(_08062_),
    .Y(_08103_));
 o21ai_1 _12700_ (.A1(_07080_),
    .A2(\digitop_pav2.access_inst.access_check0.fg_i[9] ),
    .B1(_07073_),
    .Y(_08104_));
 a21oi_2 _12701_ (.A1(net1694),
    .A2(_08033_),
    .B1(net1699),
    .Y(_08105_));
 nor2_1 _12702_ (.A(_07334_),
    .B(_08105_),
    .Y(_08106_));
 or2_1 _12703_ (.A(_07334_),
    .B(_08105_),
    .X(_08107_));
 o2111a_2 _12704_ (.A1(net1151),
    .A2(_07962_),
    .B1(net1318),
    .C1(net1065),
    .D1(net1256),
    .X(_08108_));
 a21oi_4 _12705_ (.A1(_07497_),
    .A2(net1016),
    .B1(_08108_),
    .Y(_08109_));
 a21o_1 _12706_ (.A1(_07497_),
    .A2(net1016),
    .B1(_08108_),
    .X(_08110_));
 or3_1 _12707_ (.A(net1150),
    .B(net1151),
    .C(net1016),
    .X(_08111_));
 and3b_1 _12708_ (.A_N(_07494_),
    .B(_08111_),
    .C(_07033_),
    .X(_08112_));
 or3b_2 _12709_ (.A(\digitop_pav2.access_inst.access_check0.ctrl_wcknzero_ck ),
    .B(_07494_),
    .C_N(_08111_),
    .X(_08113_));
 or3_1 _12710_ (.A(_07032_),
    .B(net1148),
    .C(net201),
    .X(_08114_));
 nor2_1 _12711_ (.A(\digitop_pav2.access_inst.access_check0.fg_i[2] ),
    .B(net195),
    .Y(_08115_));
 nand2_1 _12712_ (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[4] ),
    .B(\digitop_pav2.access_inst.access_proc0.proc_crc_check[3] ),
    .Y(_08116_));
 nand2_1 _12713_ (.A(net1036),
    .B(_08116_),
    .Y(_08117_));
 nand2_4 _12714_ (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[1] ),
    .B(_07026_),
    .Y(_08118_));
 nor2_4 _12715_ (.A(_08117_),
    .B(_08118_),
    .Y(_08119_));
 nand2_1 _12716_ (.A(net1155),
    .B(_08116_),
    .Y(_08120_));
 nor2_1 _12717_ (.A(_07476_),
    .B(_08120_),
    .Y(_08121_));
 and2_1 _12718_ (.A(net382),
    .B(_08121_),
    .X(_08122_));
 a32o_1 _12719_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[3] ),
    .A2(net382),
    .A3(_08119_),
    .B1(net342),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[3] ),
    .X(_08123_));
 and4_1 _12720_ (.A(_07025_),
    .B(net1049),
    .C(net1155),
    .D(_08116_),
    .X(_08124_));
 and2_1 _12721_ (.A(net384),
    .B(_08124_),
    .X(_08125_));
 nor2_2 _12722_ (.A(_08118_),
    .B(_08120_),
    .Y(_08126_));
 and2_2 _12723_ (.A(net383),
    .B(_08126_),
    .X(_08127_));
 a221o_1 _12724_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[3] ),
    .A2(net341),
    .B1(_08127_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[3] ),
    .C1(_08123_),
    .X(_08128_));
 and2_2 _12725_ (.A(_07478_),
    .B(_08116_),
    .X(_08129_));
 nand2_1 _12726_ (.A(_07478_),
    .B(_08116_),
    .Y(_08130_));
 nand2_1 _12727_ (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[1] ),
    .B(net1049),
    .Y(_08131_));
 nor2_1 _12728_ (.A(_08120_),
    .B(_08131_),
    .Y(_08132_));
 a31o_1 _12729_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[3] ),
    .A2(net382),
    .A3(net977),
    .B1(net979),
    .X(_08133_));
 nor3_1 _12730_ (.A(net366),
    .B(_08117_),
    .C(_08131_),
    .Y(_08134_));
 and4_1 _12731_ (.A(_07025_),
    .B(net1049),
    .C(net1036),
    .D(_08116_),
    .X(_08135_));
 and2_1 _12732_ (.A(net384),
    .B(_08135_),
    .X(_08136_));
 a221o_1 _12733_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[3] ),
    .A2(net339),
    .B1(net338),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[3] ),
    .C1(_08133_),
    .X(_08137_));
 nand2_1 _12734_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[3] ),
    .B(net387),
    .Y(_08138_));
 o2bb2a_1 _12735_ (.A1_N(net979),
    .A2_N(_08138_),
    .B1(_08137_),
    .B2(_08128_),
    .X(_08139_));
 xnor2_1 _12736_ (.A(net1126),
    .B(_08139_),
    .Y(_08140_));
 nand2_2 _12737_ (.A(_07032_),
    .B(_07564_),
    .Y(_08141_));
 and2_1 _12738_ (.A(net1068),
    .B(_08141_),
    .X(_08142_));
 nand2_1 _12739_ (.A(net1068),
    .B(_08141_),
    .Y(_08143_));
 nand2_1 _12740_ (.A(net1149),
    .B(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[3] ),
    .Y(_08144_));
 o211a_1 _12741_ (.A1(net1149),
    .A2(_08140_),
    .B1(_08144_),
    .C1(net196),
    .X(_08145_));
 o32a_1 _12742_ (.A1(_08115_),
    .A2(_08143_),
    .A3(_08145_),
    .B1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[3] ),
    .B2(net1068),
    .X(_08146_));
 and3_2 _12743_ (.A(net818),
    .B(net1016),
    .C(_08035_),
    .X(_08147_));
 and4_4 _12744_ (.A(net1081),
    .B(net1075),
    .C(_07531_),
    .D(_07535_),
    .X(_08148_));
 mux2_1 _12745_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[3] ),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[2] ),
    .S(_08148_),
    .X(_08149_));
 a21oi_1 _12746_ (.A1(_08147_),
    .A2(_08149_),
    .B1(net959),
    .Y(_08150_));
 a211o_1 _12747_ (.A1(net959),
    .A2(_08146_),
    .B1(_08150_),
    .C1(net961),
    .X(_08151_));
 a21oi_1 _12748_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[2] ),
    .A2(net961),
    .B1(net805),
    .Y(_08152_));
 o2bb2a_2 _12749_ (.A1_N(_08152_),
    .A2_N(_08151_),
    .B1(net803),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[3] ),
    .X(_08153_));
 and2_1 _12750_ (.A(net195),
    .B(_08141_),
    .X(_08154_));
 nand2_1 _12751_ (.A(net195),
    .B(_08141_),
    .Y(_08155_));
 and3_1 _12752_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[4] ),
    .B(net376),
    .C(_08119_),
    .X(_08156_));
 a221o_1 _12753_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[4] ),
    .A2(_08127_),
    .B1(net340),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[4] ),
    .C1(_08156_),
    .X(_08157_));
 a32o_1 _12754_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[4] ),
    .A2(net376),
    .A3(net977),
    .B1(net342),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[4] ),
    .X(_08158_));
 a221o_1 _12755_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[4] ),
    .A2(net341),
    .B1(_08136_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[4] ),
    .C1(_08158_),
    .X(_08159_));
 and2_1 _12756_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[4] ),
    .B(net376),
    .X(_08160_));
 a311o_1 _12757_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[4] ),
    .A2(net376),
    .A3(net979),
    .B1(_08157_),
    .C1(_08159_),
    .X(_08161_));
 nor2_1 _12758_ (.A(net1123),
    .B(_08161_),
    .Y(_08162_));
 a21o_1 _12759_ (.A1(net1123),
    .A2(_08161_),
    .B1(net1146),
    .X(_08163_));
 a2bb2o_1 _12760_ (.A1_N(_08162_),
    .A2_N(_08163_),
    .B1(net1146),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[4] ),
    .X(_08164_));
 o22a_1 _12761_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[3] ),
    .A2(net195),
    .B1(net193),
    .B2(_08164_),
    .X(_08165_));
 a2bb2o_1 _12762_ (.A1_N(net1070),
    .A2_N(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[4] ),
    .B1(_08142_),
    .B2(_08165_),
    .X(_08166_));
 mux2_1 _12763_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[4] ),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[3] ),
    .S(_08148_),
    .X(_08167_));
 a21o_1 _12764_ (.A1(_08147_),
    .A2(_08167_),
    .B1(net959),
    .X(_08168_));
 o211a_1 _12765_ (.A1(net958),
    .A2(_08166_),
    .B1(_08168_),
    .C1(_08109_),
    .X(_08169_));
 a21o_1 _12766_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[3] ),
    .A2(net960),
    .B1(net804),
    .X(_08170_));
 o22a_2 _12767_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[4] ),
    .A2(net803),
    .B1(_08169_),
    .B2(_08170_),
    .X(_08171_));
 and2_1 _12768_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[9] ),
    .B(net367),
    .X(_08172_));
 and2_1 _12769_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[9] ),
    .B(net368),
    .X(_08173_));
 a32o_1 _12770_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[9] ),
    .A2(net367),
    .A3(_08119_),
    .B1(net339),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[9] ),
    .X(_08174_));
 a221o_1 _12771_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[9] ),
    .A2(net341),
    .B1(net976),
    .B2(_08172_),
    .C1(_08174_),
    .X(_08175_));
 a32o_1 _12772_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[9] ),
    .A2(net367),
    .A3(_08135_),
    .B1(net342),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[9] ),
    .X(_08176_));
 a211o_1 _12773_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[9] ),
    .A2(_08127_),
    .B1(net978),
    .C1(_08176_),
    .X(_08177_));
 and2_1 _12774_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[9] ),
    .B(net371),
    .X(_08178_));
 o22a_1 _12775_ (.A1(_08175_),
    .A2(_08177_),
    .B1(_08178_),
    .B2(_08129_),
    .X(_08179_));
 xor2_1 _12776_ (.A(net1106),
    .B(_08179_),
    .X(_08180_));
 mux2_1 _12777_ (.A0(_08180_),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[9] ),
    .S(net1146),
    .X(_08181_));
 o22a_1 _12778_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[8] ),
    .A2(net195),
    .B1(net193),
    .B2(_08181_),
    .X(_08182_));
 a2bb2o_1 _12779_ (.A1_N(net1070),
    .A2_N(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[9] ),
    .B1(_08142_),
    .B2(_08182_),
    .X(_08183_));
 mux2_1 _12780_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[9] ),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[8] ),
    .S(_08148_),
    .X(_08184_));
 a21o_1 _12781_ (.A1(_08147_),
    .A2(_08184_),
    .B1(net959),
    .X(_08185_));
 o211a_1 _12782_ (.A1(net958),
    .A2(_08183_),
    .B1(_08185_),
    .C1(_08109_),
    .X(_08186_));
 a21o_1 _12783_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[8] ),
    .A2(net960),
    .B1(net804),
    .X(_08187_));
 o22a_2 _12784_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[9] ),
    .A2(net803),
    .B1(_08186_),
    .B2(_08187_),
    .X(_08188_));
 and2_2 _12785_ (.A(net383),
    .B(_08119_),
    .X(_08189_));
 and2_1 _12786_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[13] ),
    .B(net373),
    .X(_08190_));
 and3_1 _12787_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[13] ),
    .B(net375),
    .C(net976),
    .X(_08191_));
 a31o_1 _12788_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[13] ),
    .A2(net375),
    .A3(_08126_),
    .B1(_08191_),
    .X(_08192_));
 a221o_1 _12789_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[13] ),
    .A2(net338),
    .B1(_08189_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[13] ),
    .C1(_08192_),
    .X(_08193_));
 a31o_1 _12790_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[13] ),
    .A2(net376),
    .A3(_08124_),
    .B1(net979),
    .X(_08194_));
 a221o_1 _12791_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[13] ),
    .A2(net342),
    .B1(net339),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[13] ),
    .C1(_08194_),
    .X(_08195_));
 and2_1 _12792_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[13] ),
    .B(net376),
    .X(_08196_));
 o22a_1 _12793_ (.A1(_08193_),
    .A2(_08195_),
    .B1(_08196_),
    .B2(_08129_),
    .X(_08197_));
 xnor2_1 _12794_ (.A(net1093),
    .B(_08197_),
    .Y(_08198_));
 mux2_1 _12795_ (.A0(_08198_),
    .A1(_07103_),
    .S(net1147),
    .X(_08199_));
 o221a_1 _12796_ (.A1(net1319),
    .A2(net195),
    .B1(net193),
    .B2(_08199_),
    .C1(net1068),
    .X(_08200_));
 a211o_1 _12797_ (.A1(net1039),
    .A2(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[13] ),
    .B1(net958),
    .C1(_08200_),
    .X(_08201_));
 and2_2 _12798_ (.A(net958),
    .B(_08147_),
    .X(_08202_));
 mux2_1 _12799_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[13] ),
    .A1(net1318),
    .S(_08148_),
    .X(_08203_));
 nand2_1 _12800_ (.A(_08202_),
    .B(_08203_),
    .Y(_08204_));
 and3_1 _12801_ (.A(_08109_),
    .B(_08201_),
    .C(_08204_),
    .X(_08205_));
 a31o_1 _12802_ (.A1(net1319),
    .A2(_07497_),
    .A3(net1016),
    .B1(net805),
    .X(_08206_));
 a2bb2o_2 _12803_ (.A1_N(_08205_),
    .A2_N(_08206_),
    .B1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[13] ),
    .B2(net805),
    .X(_08207_));
 and2_1 _12804_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[6] ),
    .B(net380),
    .X(_08208_));
 a22o_1 _12805_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[6] ),
    .A2(net341),
    .B1(_08189_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[6] ),
    .X(_08209_));
 a211o_1 _12806_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[6] ),
    .A2(net340),
    .B1(_08209_),
    .C1(net979),
    .X(_08210_));
 a32o_1 _12807_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[6] ),
    .A2(net381),
    .A3(_08126_),
    .B1(net342),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[6] ),
    .X(_08211_));
 a32o_1 _12808_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[6] ),
    .A2(net383),
    .A3(net977),
    .B1(_08136_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[6] ),
    .X(_08212_));
 and2_1 _12809_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[6] ),
    .B(net385),
    .X(_08213_));
 o32a_1 _12810_ (.A1(_08210_),
    .A2(_08211_),
    .A3(_08212_),
    .B1(_08213_),
    .B2(_08129_),
    .X(_08214_));
 nand2_1 _12811_ (.A(net1117),
    .B(_08214_),
    .Y(_08215_));
 o21ba_1 _12812_ (.A1(net1117),
    .A2(_08214_),
    .B1_N(net1146),
    .X(_08216_));
 a22o_1 _12813_ (.A1(net1146),
    .A2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[6] ),
    .B1(_08215_),
    .B2(_08216_),
    .X(_08217_));
 a31o_1 _12814_ (.A1(net1066),
    .A2(\digitop_pav2.access_inst.access_check0.fg_i[5] ),
    .A3(net193),
    .B1(net1038),
    .X(_08218_));
 a21oi_1 _12815_ (.A1(_08154_),
    .A2(_08217_),
    .B1(_08218_),
    .Y(_08219_));
 a211oi_1 _12816_ (.A1(net1038),
    .A2(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[6] ),
    .B1(net958),
    .C1(_08219_),
    .Y(_08220_));
 or4bb_4 _12817_ (.A(_07532_),
    .B(net1081),
    .C_N(net1075),
    .D_N(_07535_),
    .X(_08221_));
 mux2_1 _12818_ (.A0(\digitop_pav2.access_inst.access_check0.fg_i[5] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[6] ),
    .S(_08221_),
    .X(_08222_));
 a211o_1 _12819_ (.A1(_08202_),
    .A2(_08222_),
    .B1(_08220_),
    .C1(net960),
    .X(_08223_));
 a21oi_1 _12820_ (.A1(_07097_),
    .A2(net960),
    .B1(net804),
    .Y(_08224_));
 a22o_2 _12821_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[6] ),
    .A2(net804),
    .B1(_08223_),
    .B2(_08224_),
    .X(_08225_));
 a21o_1 _12822_ (.A1(_07497_),
    .A2(net1016),
    .B1(net805),
    .X(_08226_));
 inv_2 _12823_ (.A(_08226_),
    .Y(_08227_));
 nand2_1 _12824_ (.A(net1068),
    .B(net195),
    .Y(_08228_));
 and3_1 _12825_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[15] ),
    .B(net368),
    .C(net976),
    .X(_08229_));
 a32o_1 _12826_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[15] ),
    .A2(net367),
    .A3(_08119_),
    .B1(net338),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[15] ),
    .X(_08230_));
 a31o_1 _12827_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[15] ),
    .A2(net367),
    .A3(_08126_),
    .B1(_08229_),
    .X(_08231_));
 a211o_1 _12828_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[15] ),
    .A2(net339),
    .B1(_08231_),
    .C1(net978),
    .X(_08232_));
 a221o_1 _12829_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[15] ),
    .A2(net342),
    .B1(net341),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[15] ),
    .C1(_08232_),
    .X(_08233_));
 nand2_1 _12830_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[15] ),
    .B(net372),
    .Y(_08234_));
 o2bb2a_1 _12831_ (.A1_N(net978),
    .A2_N(_08234_),
    .B1(_08233_),
    .B2(_08230_),
    .X(_08235_));
 xnor2_1 _12832_ (.A(_07061_),
    .B(_08235_),
    .Y(_08236_));
 mux2_1 _12833_ (.A0(_08236_),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[15] ),
    .S(net1149),
    .X(_08237_));
 a21o_1 _12834_ (.A1(_08141_),
    .A2(_08237_),
    .B1(_08228_),
    .X(_08238_));
 nand2_1 _12835_ (.A(net1039),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[15] ),
    .Y(_08239_));
 a31o_1 _12836_ (.A1(_08112_),
    .A2(_08238_),
    .A3(_08239_),
    .B1(_08108_),
    .X(_08240_));
 a22o_2 _12837_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[15] ),
    .A2(net805),
    .B1(_08227_),
    .B2(_08240_),
    .X(_08241_));
 xnor2_1 _12838_ (.A(_08050_),
    .B(_08241_),
    .Y(_08242_));
 nor2_1 _12839_ (.A(\digitop_pav2.access_inst.access_check0.fg_i[1] ),
    .B(net196),
    .Y(_08243_));
 and3_1 _12840_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[2] ),
    .B(net376),
    .C(_08126_),
    .X(_08244_));
 a221o_1 _12841_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[2] ),
    .A2(net341),
    .B1(net340),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[2] ),
    .C1(_08244_),
    .X(_08245_));
 and2_1 _12842_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[2] ),
    .B(net375),
    .X(_08246_));
 a32o_1 _12843_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[2] ),
    .A2(net381),
    .A3(net976),
    .B1(_08189_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[2] ),
    .X(_08247_));
 a221o_1 _12844_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[2] ),
    .A2(_08136_),
    .B1(_08246_),
    .B2(_08121_),
    .C1(_08247_),
    .X(_08248_));
 a311o_1 _12845_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ),
    .A2(net376),
    .A3(net979),
    .B1(_08245_),
    .C1(_08248_),
    .X(_08249_));
 nor2_1 _12846_ (.A(net1127),
    .B(_08249_),
    .Y(_08250_));
 and2_1 _12847_ (.A(net1127),
    .B(_08249_),
    .X(_08251_));
 nand2_1 _12848_ (.A(net1149),
    .B(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[2] ),
    .Y(_08252_));
 o311a_1 _12849_ (.A1(net1149),
    .A2(_08250_),
    .A3(_08251_),
    .B1(_08252_),
    .C1(net196),
    .X(_08253_));
 o32a_1 _12850_ (.A1(_08143_),
    .A2(_08243_),
    .A3(_08253_),
    .B1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[2] ),
    .B2(net1068),
    .X(_08254_));
 mux2_1 _12851_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[2] ),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[1] ),
    .S(_08148_),
    .X(_08255_));
 a21oi_1 _12852_ (.A1(_08147_),
    .A2(_08255_),
    .B1(net959),
    .Y(_08256_));
 a211o_1 _12853_ (.A1(net959),
    .A2(_08254_),
    .B1(_08256_),
    .C1(net961),
    .X(_08257_));
 a21oi_1 _12854_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[1] ),
    .A2(net961),
    .B1(net804),
    .Y(_08258_));
 o2bb2a_1 _12855_ (.A1_N(_08258_),
    .A2_N(_08257_),
    .B1(net803),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[2] ),
    .X(_08259_));
 and3_1 _12856_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[10] ),
    .B(net375),
    .C(_08124_),
    .X(_08260_));
 a31o_1 _12857_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[10] ),
    .A2(net375),
    .A3(net976),
    .B1(_08260_),
    .X(_08261_));
 a221o_1 _12858_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ),
    .A2(_08122_),
    .B1(_08127_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ),
    .C1(_08261_),
    .X(_08262_));
 a31o_1 _12859_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[10] ),
    .A2(net375),
    .A3(_08119_),
    .B1(net979),
    .X(_08263_));
 a221o_1 _12860_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[10] ),
    .A2(net339),
    .B1(net338),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[10] ),
    .C1(_08263_),
    .X(_08264_));
 nand2_1 _12861_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[10] ),
    .B(net385),
    .Y(_08265_));
 o2bb2a_1 _12862_ (.A1_N(net979),
    .A2_N(_08265_),
    .B1(_08264_),
    .B2(_08262_),
    .X(_08266_));
 or2_1 _12863_ (.A(net1102),
    .B(_08266_),
    .X(_08267_));
 a21oi_1 _12864_ (.A1(net1102),
    .A2(_08266_),
    .B1(net1146),
    .Y(_08268_));
 a22o_1 _12865_ (.A1(net1146),
    .A2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[10] ),
    .B1(_08267_),
    .B2(_08268_),
    .X(_08269_));
 o22a_1 _12866_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[9] ),
    .A2(net195),
    .B1(net193),
    .B2(_08269_),
    .X(_08270_));
 a2bb2o_1 _12867_ (.A1_N(net1068),
    .A2_N(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[10] ),
    .B1(_08142_),
    .B2(_08270_),
    .X(_08271_));
 mux2_1 _12868_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[10] ),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[9] ),
    .S(_08148_),
    .X(_08272_));
 a21o_1 _12869_ (.A1(_08147_),
    .A2(_08272_),
    .B1(net959),
    .X(_08273_));
 o211a_1 _12870_ (.A1(net958),
    .A2(_08271_),
    .B1(_08273_),
    .C1(_08109_),
    .X(_08274_));
 a21o_1 _12871_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[9] ),
    .A2(net960),
    .B1(net804),
    .X(_08275_));
 o22a_2 _12872_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[10] ),
    .A2(net803),
    .B1(_08274_),
    .B2(_08275_),
    .X(_08276_));
 xnor2_1 _12873_ (.A(_08075_),
    .B(_08276_),
    .Y(_08277_));
 a32o_1 _12874_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[1] ),
    .A2(net382),
    .A3(_08126_),
    .B1(_08189_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[1] ),
    .X(_08278_));
 and2_1 _12875_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[1] ),
    .B(net382),
    .X(_08279_));
 a32o_1 _12876_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[1] ),
    .A2(net383),
    .A3(net977),
    .B1(_08125_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[1] ),
    .X(_08280_));
 a221o_1 _12877_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[1] ),
    .A2(_08122_),
    .B1(_08135_),
    .B2(_08279_),
    .C1(_08278_),
    .X(_08281_));
 a211o_1 _12878_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[1] ),
    .A2(net340),
    .B1(_08280_),
    .C1(net979),
    .X(_08282_));
 a21o_1 _12879_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[1] ),
    .A2(net383),
    .B1(_08129_),
    .X(_08283_));
 o21ai_1 _12880_ (.A1(_08281_),
    .A2(_08282_),
    .B1(_08283_),
    .Y(_08284_));
 xnor2_1 _12881_ (.A(net1132),
    .B(_08284_),
    .Y(_08285_));
 mux2_1 _12882_ (.A0(_08285_),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[1] ),
    .S(net1147),
    .X(_08286_));
 o22a_1 _12883_ (.A1(net1324),
    .A2(net195),
    .B1(net193),
    .B2(_08286_),
    .X(_08287_));
 a2bb2o_1 _12884_ (.A1_N(net1068),
    .A2_N(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[1] ),
    .B1(_08142_),
    .B2(_08287_),
    .X(_08288_));
 mux2_1 _12885_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[1] ),
    .A1(net1324),
    .S(_08148_),
    .X(_08289_));
 a21o_1 _12886_ (.A1(_08147_),
    .A2(_08289_),
    .B1(net959),
    .X(_08290_));
 o211a_1 _12887_ (.A1(net958),
    .A2(_08288_),
    .B1(_08290_),
    .C1(_08109_),
    .X(_08291_));
 a21o_1 _12888_ (.A1(net1324),
    .A2(net961),
    .B1(net805),
    .X(_08292_));
 o22a_2 _12889_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[1] ),
    .A2(net803),
    .B1(_08291_),
    .B2(_08292_),
    .X(_08293_));
 a32o_1 _12890_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[12] ),
    .A2(net367),
    .A3(_08126_),
    .B1(net342),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[12] ),
    .X(_08294_));
 a221o_1 _12891_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[12] ),
    .A2(net338),
    .B1(_08189_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[12] ),
    .C1(_08294_),
    .X(_08295_));
 a32o_1 _12892_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[12] ),
    .A2(net376),
    .A3(net976),
    .B1(net341),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[12] ),
    .X(_08296_));
 a211o_1 _12893_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[12] ),
    .A2(net339),
    .B1(_08296_),
    .C1(net978),
    .X(_08297_));
 nand2_1 _12894_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[12] ),
    .B(net370),
    .Y(_08298_));
 o2bb2a_1 _12895_ (.A1_N(net978),
    .A2_N(_08298_),
    .B1(_08297_),
    .B2(_08295_),
    .X(_08299_));
 xnor2_1 _12896_ (.A(net1035),
    .B(_08299_),
    .Y(_08300_));
 mux2_1 _12897_ (.A0(_08300_),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[12] ),
    .S(net1149),
    .X(_08301_));
 a31o_1 _12898_ (.A1(net1066),
    .A2(\digitop_pav2.access_inst.access_check0.fg_i[11] ),
    .A3(net193),
    .B1(net1038),
    .X(_08302_));
 a21oi_1 _12899_ (.A1(_08154_),
    .A2(_08301_),
    .B1(_08302_),
    .Y(_08303_));
 a211oi_1 _12900_ (.A1(net1039),
    .A2(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[12] ),
    .B1(_08113_),
    .C1(_08303_),
    .Y(_08304_));
 mux2_1 _12901_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[12] ),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[11] ),
    .S(_08148_),
    .X(_08305_));
 a211o_1 _12902_ (.A1(_08202_),
    .A2(_08305_),
    .B1(_08304_),
    .C1(net961),
    .X(_08306_));
 o21a_1 _12903_ (.A1(net1790),
    .A2(_08109_),
    .B1(net803),
    .X(_08307_));
 a22o_2 _12904_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[12] ),
    .A2(net805),
    .B1(_08306_),
    .B2(_08307_),
    .X(_08308_));
 nand2_1 _12905_ (.A(\digitop_pav2.access_inst.acc_wcknzero_o ),
    .B(_08108_),
    .Y(_08309_));
 and3_1 _12906_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[0] ),
    .B(net382),
    .C(_08124_),
    .X(_08310_));
 and2_1 _12907_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[0] ),
    .B(net382),
    .X(_08311_));
 a31o_1 _12908_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[0] ),
    .A2(net382),
    .A3(_08119_),
    .B1(_08310_),
    .X(_08312_));
 a31o_1 _12909_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[0] ),
    .A2(net382),
    .A3(net977),
    .B1(_08130_),
    .X(_08313_));
 a22o_1 _12910_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ),
    .A2(_08122_),
    .B1(_08127_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[0] ),
    .X(_08314_));
 a221o_1 _12911_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[0] ),
    .A2(net340),
    .B1(_08135_),
    .B2(_08311_),
    .C1(_08314_),
    .X(_08315_));
 a21o_1 _12912_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[0] ),
    .A2(net383),
    .B1(_08129_),
    .X(_08316_));
 o31a_1 _12913_ (.A1(_08312_),
    .A2(_08313_),
    .A3(_08315_),
    .B1(_08316_),
    .X(_08317_));
 xnor2_1 _12914_ (.A(net1135),
    .B(_08317_),
    .Y(_08318_));
 nand2_1 _12915_ (.A(net1149),
    .B(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[0] ),
    .Y(_08319_));
 o211ai_1 _12916_ (.A1(net1149),
    .A2(_08318_),
    .B1(_08319_),
    .C1(net196),
    .Y(_08320_));
 o211ai_1 _12917_ (.A1(\digitop_pav2.access_inst.acc_wcknzero_o ),
    .A2(net196),
    .B1(_08141_),
    .C1(_08320_),
    .Y(_08321_));
 mux2_1 _12918_ (.A0(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[0] ),
    .A1(_08321_),
    .S(net1070),
    .X(_08322_));
 o31a_1 _12919_ (.A1(_08108_),
    .A2(_08113_),
    .A3(_08322_),
    .B1(_08309_),
    .X(_08323_));
 o2bb2a_2 _12920_ (.A1_N(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[0] ),
    .A2_N(net805),
    .B1(_08226_),
    .B2(_08323_),
    .X(_08324_));
 xnor2_1 _12921_ (.A(_08060_),
    .B(_08324_),
    .Y(_08325_));
 and3_1 _12922_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ),
    .B(net375),
    .C(_08124_),
    .X(_08326_));
 a32o_1 _12923_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[7] ),
    .A2(net375),
    .A3(net976),
    .B1(net339),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[7] ),
    .X(_08327_));
 a311o_1 _12924_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ),
    .A2(net375),
    .A3(_08121_),
    .B1(_08326_),
    .C1(_08327_),
    .X(_08328_));
 a31o_1 _12925_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[7] ),
    .A2(net367),
    .A3(_08119_),
    .B1(net978),
    .X(_08329_));
 a221o_1 _12926_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[7] ),
    .A2(_08127_),
    .B1(net338),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ),
    .C1(_08329_),
    .X(_08330_));
 and2_1 _12927_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ),
    .B(net371),
    .X(_08331_));
 o22a_1 _12928_ (.A1(_08328_),
    .A2(_08330_),
    .B1(_08331_),
    .B2(_08129_),
    .X(_08332_));
 xor2_1 _12929_ (.A(net1114),
    .B(_08332_),
    .X(_08333_));
 mux2_1 _12930_ (.A0(_08333_),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[7] ),
    .S(net1147),
    .X(_08334_));
 o22a_1 _12931_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[6] ),
    .A2(net195),
    .B1(net193),
    .B2(_08334_),
    .X(_08335_));
 o2bb2a_1 _12932_ (.A1_N(_08142_),
    .A2_N(_08335_),
    .B1(net1068),
    .B2(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[7] ),
    .X(_08336_));
 mux2_1 _12933_ (.A0(\digitop_pav2.access_inst.access_check0.fg_i[6] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[7] ),
    .S(_08221_),
    .X(_08337_));
 a21o_1 _12934_ (.A1(_08147_),
    .A2(_08337_),
    .B1(net959),
    .X(_08338_));
 a21oi_1 _12935_ (.A1(net959),
    .A2(_08336_),
    .B1(net960),
    .Y(_08339_));
 a221o_1 _12936_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[6] ),
    .A2(net960),
    .B1(_08338_),
    .B2(_08339_),
    .C1(net804),
    .X(_08340_));
 o21ai_2 _12937_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[7] ),
    .A2(net803),
    .B1(_08340_),
    .Y(_08341_));
 a32o_1 _12938_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[8] ),
    .A2(net368),
    .A3(_08126_),
    .B1(net341),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[8] ),
    .X(_08342_));
 a221o_1 _12939_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[8] ),
    .A2(net342),
    .B1(net339),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[8] ),
    .C1(_08342_),
    .X(_08343_));
 a32o_1 _12940_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[8] ),
    .A2(net368),
    .A3(net976),
    .B1(net338),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[8] ),
    .X(_08344_));
 a211o_1 _12941_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[8] ),
    .A2(_08189_),
    .B1(_08344_),
    .C1(net978),
    .X(_08345_));
 nand2_1 _12942_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[8] ),
    .B(net374),
    .Y(_08346_));
 o2bb2a_1 _12943_ (.A1_N(net978),
    .A2_N(_08346_),
    .B1(_08345_),
    .B2(_08343_),
    .X(_08347_));
 xnor2_2 _12944_ (.A(_07079_),
    .B(_08347_),
    .Y(_08348_));
 mux2_1 _12945_ (.A0(_08348_),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[8] ),
    .S(net1146),
    .X(_08349_));
 a31o_1 _12946_ (.A1(net1066),
    .A2(\digitop_pav2.access_inst.access_check0.fg_i[7] ),
    .A3(net193),
    .B1(net1038),
    .X(_08350_));
 a21oi_1 _12947_ (.A1(_08154_),
    .A2(_08349_),
    .B1(_08350_),
    .Y(_08351_));
 a211oi_1 _12948_ (.A1(net1039),
    .A2(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[8] ),
    .B1(net958),
    .C1(_08351_),
    .Y(_08352_));
 mux2_1 _12949_ (.A0(\digitop_pav2.access_inst.access_check0.fg_i[7] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[8] ),
    .S(_08221_),
    .X(_08353_));
 a211o_1 _12950_ (.A1(_08202_),
    .A2(_08353_),
    .B1(_08352_),
    .C1(net960),
    .X(_08354_));
 a21oi_1 _12951_ (.A1(_07099_),
    .A2(net960),
    .B1(net804),
    .Y(_08355_));
 a22o_1 _12952_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[8] ),
    .A2(net804),
    .B1(_08354_),
    .B2(_08355_),
    .X(_08356_));
 and3_1 _12953_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[5] ),
    .B(net382),
    .C(_08119_),
    .X(_08357_));
 a221o_1 _12954_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[5] ),
    .A2(_08127_),
    .B1(net340),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[5] ),
    .C1(_08357_),
    .X(_08358_));
 and2_1 _12955_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[5] ),
    .B(net383),
    .X(_08359_));
 a32o_1 _12956_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[5] ),
    .A2(net383),
    .A3(net977),
    .B1(_08359_),
    .B2(_08121_),
    .X(_08360_));
 a221o_1 _12957_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[5] ),
    .A2(_08125_),
    .B1(net338),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[5] ),
    .C1(_08360_),
    .X(_08361_));
 a311o_1 _12958_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[5] ),
    .A2(net383),
    .A3(_08130_),
    .B1(_08358_),
    .C1(_08361_),
    .X(_08362_));
 nand2_1 _12959_ (.A(net1120),
    .B(_08362_),
    .Y(_08363_));
 o21ba_1 _12960_ (.A1(net1120),
    .A2(_08362_),
    .B1_N(net1146),
    .X(_08364_));
 a22o_1 _12961_ (.A1(net1146),
    .A2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[5] ),
    .B1(_08363_),
    .B2(_08364_),
    .X(_08365_));
 a31o_1 _12962_ (.A1(net1066),
    .A2(net1323),
    .A3(_08155_),
    .B1(net1038),
    .X(_08366_));
 a21oi_1 _12963_ (.A1(_08154_),
    .A2(_08365_),
    .B1(_08366_),
    .Y(_08367_));
 a211oi_1 _12964_ (.A1(net1039),
    .A2(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[5] ),
    .B1(net958),
    .C1(_08367_),
    .Y(_08368_));
 mux2_1 _12965_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[5] ),
    .A1(net1323),
    .S(_08148_),
    .X(_08369_));
 a211o_1 _12966_ (.A1(_08202_),
    .A2(_08369_),
    .B1(_08368_),
    .C1(net960),
    .X(_08370_));
 o21a_1 _12967_ (.A1(net1323),
    .A2(_08109_),
    .B1(net803),
    .X(_08371_));
 a22o_1 _12968_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[5] ),
    .A2(net804),
    .B1(_08370_),
    .B2(_08371_),
    .X(_08372_));
 a22o_1 _12969_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[11] ),
    .A2(net341),
    .B1(net339),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[11] ),
    .X(_08373_));
 a31o_1 _12970_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[11] ),
    .A2(net368),
    .A3(net976),
    .B1(net978),
    .X(_08374_));
 a22o_1 _12971_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[11] ),
    .A2(net338),
    .B1(_08189_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[11] ),
    .X(_08375_));
 a221o_1 _12972_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[11] ),
    .A2(net342),
    .B1(_08127_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[11] ),
    .C1(_08375_),
    .X(_08376_));
 and2_1 _12973_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[11] ),
    .B(net372),
    .X(_08377_));
 o32a_1 _12974_ (.A1(_08373_),
    .A2(_08374_),
    .A3(_08376_),
    .B1(_08377_),
    .B2(_08129_),
    .X(_08378_));
 xor2_1 _12975_ (.A(net1098),
    .B(_08378_),
    .X(_08379_));
 mux2_1 _12976_ (.A0(_08379_),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[11] ),
    .S(net1147),
    .X(_08380_));
 a31o_1 _12977_ (.A1(net1066),
    .A2(\digitop_pav2.access_inst.access_check0.fg_i[10] ),
    .A3(net193),
    .B1(net1038),
    .X(_08381_));
 a21oi_1 _12978_ (.A1(_08154_),
    .A2(_08380_),
    .B1(_08381_),
    .Y(_08382_));
 a211oi_1 _12979_ (.A1(net1039),
    .A2(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[11] ),
    .B1(net958),
    .C1(_08382_),
    .Y(_08383_));
 mux2_1 _12980_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[11] ),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[10] ),
    .S(_08148_),
    .X(_08384_));
 a211o_1 _12981_ (.A1(_08202_),
    .A2(_08384_),
    .B1(_08383_),
    .C1(net961),
    .X(_08385_));
 o21a_1 _12982_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[10] ),
    .A2(_08109_),
    .B1(_08107_),
    .X(_08386_));
 a22o_1 _12983_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[11] ),
    .A2(net805),
    .B1(_08385_),
    .B2(_08386_),
    .X(_08387_));
 and2_1 _12984_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[14] ),
    .B(net367),
    .X(_08388_));
 a32o_1 _12985_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[14] ),
    .A2(net367),
    .A3(_08126_),
    .B1(net342),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[14] ),
    .X(_08389_));
 a32o_1 _12986_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[14] ),
    .A2(net375),
    .A3(net976),
    .B1(_08388_),
    .B2(_08119_),
    .X(_08390_));
 a211o_1 _12987_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[14] ),
    .A2(net338),
    .B1(_08390_),
    .C1(net978),
    .X(_08391_));
 a221o_1 _12988_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[14] ),
    .A2(net341),
    .B1(net339),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[14] ),
    .C1(_08391_),
    .X(_08392_));
 and2_1 _12989_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[14] ),
    .B(net367),
    .X(_08393_));
 o22a_1 _12990_ (.A1(_08389_),
    .A2(_08392_),
    .B1(_08393_),
    .B2(_08129_),
    .X(_08394_));
 xnor2_1 _12991_ (.A(_07083_),
    .B(_08394_),
    .Y(_08395_));
 mux2_1 _12992_ (.A0(_08395_),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[14] ),
    .S(net1147),
    .X(_08396_));
 a21oi_1 _12993_ (.A1(_08141_),
    .A2(_08396_),
    .B1(_08228_),
    .Y(_08397_));
 a2111o_1 _12994_ (.A1(net1039),
    .A2(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[14] ),
    .B1(_08108_),
    .C1(_08113_),
    .D1(_08397_),
    .X(_08398_));
 o2bb2a_2 _12995_ (.A1_N(_08227_),
    .A2_N(_08398_),
    .B1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[14] ),
    .B2(net803),
    .X(_08399_));
 xnor2_1 _12996_ (.A(_08084_),
    .B(_08399_),
    .Y(_08400_));
 xnor2_1 _12997_ (.A(_08070_),
    .B(_08356_),
    .Y(_08401_));
 a2bb2o_1 _12998_ (.A1_N(_08059_),
    .A2_N(_08259_),
    .B1(_08308_),
    .B2(_08067_),
    .X(_08402_));
 a221o_1 _12999_ (.A1(_08083_),
    .A2(_08225_),
    .B1(_08387_),
    .B2(_08064_),
    .C1(_08402_),
    .X(_08403_));
 a2bb2o_1 _13000_ (.A1_N(_08387_),
    .A2_N(_08064_),
    .B1(_08059_),
    .B2(_08259_),
    .X(_08404_));
 xnor2_1 _13001_ (.A(_08052_),
    .B(_08372_),
    .Y(_08405_));
 o221a_1 _13002_ (.A1(_08083_),
    .A2(_08225_),
    .B1(_08308_),
    .B2(_08067_),
    .C1(_08405_),
    .X(_08406_));
 or4b_1 _13003_ (.A(_08277_),
    .B(_08401_),
    .C(_08404_),
    .D_N(_08406_),
    .X(_08407_));
 a22o_1 _13004_ (.A1(_08078_),
    .A2(_08153_),
    .B1(_08171_),
    .B2(_08081_),
    .X(_08408_));
 o21ba_1 _13005_ (.A1(_08078_),
    .A2(_08153_),
    .B1_N(_08408_),
    .X(_08409_));
 o221a_1 _13006_ (.A1(_08062_),
    .A2(_08188_),
    .B1(_08293_),
    .B2(_08057_),
    .C1(_08409_),
    .X(_08410_));
 xnor2_1 _13007_ (.A(_08072_),
    .B(_08207_),
    .Y(_08411_));
 or4_1 _13008_ (.A(_08035_),
    .B(_08242_),
    .C(_08400_),
    .D(_08411_),
    .X(_08412_));
 a22o_1 _13009_ (.A1(_08057_),
    .A2(_08293_),
    .B1(_08341_),
    .B2(_08054_),
    .X(_08413_));
 a21oi_1 _13010_ (.A1(_08062_),
    .A2(_08188_),
    .B1(_08413_),
    .Y(_08414_));
 and4b_1 _13011_ (.A_N(_08412_),
    .B(_08325_),
    .C(_08410_),
    .D(_08414_),
    .X(_08415_));
 o221a_1 _13012_ (.A1(_08081_),
    .A2(_08171_),
    .B1(_08341_),
    .B2(_08054_),
    .C1(_08415_),
    .X(_08416_));
 or3b_1 _13013_ (.A(_08403_),
    .B(_08407_),
    .C_N(_08416_),
    .X(_08417_));
 a22o_1 _13014_ (.A1(_08067_),
    .A2(_08305_),
    .B1(_08384_),
    .B2(_08064_),
    .X(_08418_));
 o22ai_1 _13015_ (.A1(_08067_),
    .A2(_08305_),
    .B1(_08384_),
    .B2(_08064_),
    .Y(_08419_));
 or2_1 _13016_ (.A(_08053_),
    .B(_08369_),
    .X(_08420_));
 nand2_1 _13017_ (.A(_08053_),
    .B(_08369_),
    .Y(_08421_));
 xnor2_1 _13018_ (.A(_08055_),
    .B(_08337_),
    .Y(_08422_));
 a2bb2o_1 _13019_ (.A1_N(_08062_),
    .A2_N(_08184_),
    .B1(_08353_),
    .B2(_08070_),
    .X(_08423_));
 o2bb2a_1 _13020_ (.A1_N(_08075_),
    .A2_N(_08272_),
    .B1(_08255_),
    .B2(_08059_),
    .X(_08424_));
 o2111ai_1 _13021_ (.A1(_08075_),
    .A2(_08272_),
    .B1(_08420_),
    .C1(_08421_),
    .D1(_08424_),
    .Y(_08425_));
 o22ai_1 _13022_ (.A1(_08078_),
    .A2(_08149_),
    .B1(_08167_),
    .B2(_08081_),
    .Y(_08426_));
 a22o_1 _13023_ (.A1(_08062_),
    .A2(_08184_),
    .B1(_08289_),
    .B2(_08057_),
    .X(_08427_));
 and4_1 _13024_ (.A(_08035_),
    .B(_08050_),
    .C(_08060_),
    .D(_08084_),
    .X(_08428_));
 o221a_1 _13025_ (.A1(_08057_),
    .A2(_08289_),
    .B1(_08353_),
    .B2(_08070_),
    .C1(_08428_),
    .X(_08429_));
 or3b_1 _13026_ (.A(_08426_),
    .B(_08427_),
    .C_N(_08429_),
    .X(_08430_));
 a2bb2o_1 _13027_ (.A1_N(_08072_),
    .A2_N(_08203_),
    .B1(_08167_),
    .B2(_08081_),
    .X(_08431_));
 xnor2_1 _13028_ (.A(_08083_),
    .B(_08222_),
    .Y(_08432_));
 a22o_1 _13029_ (.A1(_08072_),
    .A2(_08203_),
    .B1(_08255_),
    .B2(_08059_),
    .X(_08433_));
 or4_1 _13030_ (.A(_08422_),
    .B(_08431_),
    .C(_08432_),
    .D(_08433_),
    .X(_08434_));
 or4_1 _13031_ (.A(_08418_),
    .B(_08419_),
    .C(_08430_),
    .D(_08434_),
    .X(_08435_));
 a2111o_1 _13032_ (.A1(_08078_),
    .A2(_08149_),
    .B1(_08423_),
    .C1(_08425_),
    .D1(_08435_),
    .X(_08436_));
 a22o_1 _13033_ (.A1(net1323),
    .A2(_08053_),
    .B1(_08057_),
    .B2(net1324),
    .X(_08437_));
 or3_1 _13034_ (.A(net1083),
    .B(_08084_),
    .C(_08104_),
    .X(_08438_));
 a221o_1 _13035_ (.A1(_07098_),
    .A2(_08054_),
    .B1(_08069_),
    .B2(_07099_),
    .C1(_08103_),
    .X(_08439_));
 o22ai_1 _13036_ (.A1(net1323),
    .A2(_08053_),
    .B1(_08057_),
    .B2(net1324),
    .Y(_08440_));
 a221o_1 _13037_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[1] ),
    .A2(_08059_),
    .B1(_08083_),
    .B2(\digitop_pav2.access_inst.access_check0.fg_i[5] ),
    .C1(_08440_),
    .X(_08441_));
 a2bb2o_1 _13038_ (.A1_N(\digitop_pav2.access_inst.access_check0.fg_i[11] ),
    .A2_N(_08067_),
    .B1(_08064_),
    .B2(\digitop_pav2.access_inst.access_check0.fg_i[10] ),
    .X(_08442_));
 a2bb2o_1 _13039_ (.A1_N(\digitop_pav2.access_inst.access_check0.fg_i[10] ),
    .A2_N(_08064_),
    .B1(_08067_),
    .B2(\digitop_pav2.access_inst.access_check0.fg_i[11] ),
    .X(_08443_));
 xnor2_1 _13040_ (.A(\digitop_pav2.access_inst.access_check0.fg_i[2] ),
    .B(_08078_),
    .Y(_08444_));
 a221o_1 _13041_ (.A1(_07095_),
    .A2(_08058_),
    .B1(_08073_),
    .B2(net1319),
    .C1(_08444_),
    .X(_08445_));
 a22o_1 _13042_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[7] ),
    .A2(_08070_),
    .B1(_08075_),
    .B2(\digitop_pav2.access_inst.access_check0.fg_i[9] ),
    .X(_08446_));
 a221o_1 _13043_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[3] ),
    .A2(_08081_),
    .B1(_08082_),
    .B2(_07097_),
    .C1(_08446_),
    .X(_08447_));
 a2111o_1 _13044_ (.A1(_07096_),
    .A2(_08080_),
    .B1(_08438_),
    .C1(_08445_),
    .D1(_08447_),
    .X(_08448_));
 a221o_1 _13045_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[6] ),
    .A2(_08055_),
    .B1(_08072_),
    .B2(net1318),
    .C1(_08437_),
    .X(_08449_));
 or4_1 _13046_ (.A(_08439_),
    .B(_08441_),
    .C(_08448_),
    .D(_08449_),
    .X(_08450_));
 or3_1 _13047_ (.A(_08442_),
    .B(_08443_),
    .C(_08450_),
    .X(_08451_));
 and4b_1 _13048_ (.A_N(net1147),
    .B(_08451_),
    .C(net1256),
    .D(\digitop_pav2.access_inst.access_check0.wr_lock_ck_i ),
    .X(_08452_));
 a311o_1 _13049_ (.A1(net1256),
    .A2(net1149),
    .A3(_08102_),
    .B1(_08452_),
    .C1(net1151),
    .X(_08453_));
 and3_1 _13050_ (.A(_08105_),
    .B(_08417_),
    .C(_08436_),
    .X(_08454_));
 and2b_1 _13051_ (.A_N(_08105_),
    .B(_08102_),
    .X(_08455_));
 o31ai_2 _13052_ (.A1(_07091_),
    .A2(_08454_),
    .A3(_08455_),
    .B1(_08453_),
    .Y(_08456_));
 a2bb2o_1 _13053_ (.A1_N(_08041_),
    .A2_N(_08456_),
    .B1(\digitop_pav2.access_inst.access_check0.write_error_reg ),
    .B2(_08040_),
    .X(_01515_));
 a31o_1 _13054_ (.A1(net1065),
    .A2(net1151),
    .A3(net1190),
    .B1(_07033_),
    .X(_08457_));
 o31ai_1 _13055_ (.A1(net1065),
    .A2(net1038),
    .A3(net1203),
    .B1(_08457_),
    .Y(_01514_));
 or2_1 _13056_ (.A(\digitop_pav2.access_inst.access_check0.mem_sign_check_sync_o ),
    .B(_07970_),
    .X(_01513_));
 a21o_1 _13057_ (.A1(net1069),
    .A2(_08038_),
    .B1(_08039_),
    .X(_01512_));
 and2_1 _13058_ (.A(\digitop_pav2.access_inst.access_check0.wr_lock_ck_i ),
    .B(_08456_),
    .X(_08458_));
 o31ai_2 _13059_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[13] ),
    .A2(\digitop_pav2.access_inst.access_check0.act_lock_st ),
    .A3(_08458_),
    .B1(net1319),
    .Y(_08459_));
 a311o_1 _13060_ (.A1(net1239),
    .A2(net811),
    .A3(_08459_),
    .B1(_07104_),
    .C1(net1206),
    .X(_08460_));
 a211o_1 _13061_ (.A1(_07604_),
    .A2(_08459_),
    .B1(net1257),
    .C1(_07321_),
    .X(_08461_));
 nor2_1 _13062_ (.A(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[2] ),
    .B(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[3] ),
    .Y(_08462_));
 or4b_1 _13063_ (.A(net1081),
    .B(net1077),
    .C(_08462_),
    .D_N(net1079),
    .X(_08463_));
 o2bb2a_1 _13064_ (.A1_N(\digitop_pav2.access_inst.access_check0.permalock_tid_i ),
    .A2_N(_07510_),
    .B1(net912),
    .B2(_08463_),
    .X(_08464_));
 o21ai_1 _13065_ (.A1(_07543_),
    .A2(_08464_),
    .B1(_08459_),
    .Y(_08465_));
 a32o_1 _13066_ (.A1(_07966_),
    .A2(_08461_),
    .A3(_08465_),
    .B1(_08460_),
    .B2(\digitop_pav2.access_inst.access_check0.lock_error_o ),
    .X(_01511_));
 nand2_1 _13067_ (.A(\digitop_pav2.access_inst.access_ctrl0.dt_acc_done_o ),
    .B(net1191),
    .Y(_08466_));
 o21ai_1 _13068_ (.A1(_07036_),
    .A2(net1191),
    .B1(_08466_),
    .Y(_01510_));
 or4_1 _13069_ (.A(\digitop_pav2.access_inst.access_ctrl0.state[1] ),
    .B(\digitop_pav2.access_inst.access_ctrl0.state[22] ),
    .C(net1205),
    .D(_07410_),
    .X(_08467_));
 nor2_1 _13070_ (.A(\digitop_pav2.access_inst.access_ctrl0.state[19] ),
    .B(_08467_),
    .Y(_08468_));
 and2b_1 _13071_ (.A_N(\digitop_pav2.access_inst.access_check0.write_error_reg ),
    .B(_08456_),
    .X(_08469_));
 or2_2 _13072_ (.A(\digitop_pav2.access_inst.access_check0.ctrl_wcknzero_ck ),
    .B(_08469_),
    .X(_08470_));
 o21ai_1 _13073_ (.A1(_07091_),
    .A2(_08470_),
    .B1(_08468_),
    .Y(_08471_));
 o22a_1 _13074_ (.A1(\digitop_pav2.access_inst.access_ctrl0.replay_nok ),
    .A2(_08468_),
    .B1(_08471_),
    .B2(\digitop_pav2.access_inst.access_ctrl0.state[5] ),
    .X(_01509_));
 and2_1 _13075_ (.A(net1240),
    .B(net1143),
    .X(_08472_));
 nor2_1 _13076_ (.A(_08467_),
    .B(_08472_),
    .Y(_08473_));
 and3_1 _13077_ (.A(net1069),
    .B(net1143),
    .C(_07575_),
    .X(_08474_));
 a21o_1 _13078_ (.A1(net1152),
    .A2(_07396_),
    .B1(_08474_),
    .X(_08475_));
 a21bo_1 _13079_ (.A1(_08470_),
    .A2(_08475_),
    .B1_N(_07554_),
    .X(_08476_));
 o31a_1 _13080_ (.A1(net1143),
    .A2(net1152),
    .A3(\digitop_pav2.access_inst.access_ctrl0.state[10] ),
    .B1(_08473_),
    .X(_08477_));
 a2bb2o_1 _13081_ (.A1_N(_07038_),
    .A2_N(_08473_),
    .B1(_08476_),
    .B2(_08477_),
    .X(_01508_));
 mux2_1 _13082_ (.A0(\digitop_pav2.access_inst.access_check0.wordcnt_i[0] ),
    .A1(net1071),
    .S(_07965_),
    .X(_01506_));
 or4b_1 _13083_ (.A(net1148),
    .B(\digitop_pav2.access_inst.access_ctrl0.state[11] ),
    .C(_07486_),
    .D_N(_08468_),
    .X(_08478_));
 mux2_1 _13084_ (.A0(net1144),
    .A1(\digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt ),
    .S(_08478_),
    .X(_01505_));
 mux2_1 _13085_ (.A0(\digitop_pav2.crc_inst.crc5_q[4] ),
    .A1(\digitop_pav2.crc_inst.crc5_q[3] ),
    .S(net1302),
    .X(_01193_));
 a21oi_1 _13086_ (.A1(\digitop_pav2.crc_inst.crc5_q[4] ),
    .A2(net1299),
    .B1(net1296),
    .Y(_08479_));
 o21ai_1 _13087_ (.A1(\digitop_pav2.crc_inst.crc5_q[4] ),
    .A2(net1299),
    .B1(_08479_),
    .Y(_08480_));
 mux2_1 _13088_ (.A0(\digitop_pav2.crc_inst.crc5_q[3] ),
    .A1(\digitop_pav2.crc_inst.crc5_q[2] ),
    .S(net1302),
    .X(_08481_));
 mux2_1 _13089_ (.A0(_07042_),
    .A1(_08481_),
    .S(_08480_),
    .X(_01192_));
 mux2_1 _13090_ (.A0(\digitop_pav2.crc_inst.crc5_q[2] ),
    .A1(\digitop_pav2.crc_inst.crc5_q[1] ),
    .S(net1302),
    .X(_01191_));
 mux2_1 _13091_ (.A0(\digitop_pav2.crc_inst.crc5_q[1] ),
    .A1(\digitop_pav2.crc_inst.crc5_q[0] ),
    .S(net1302),
    .X(_01190_));
 a21bo_1 _13092_ (.A1(net1296),
    .A2(\digitop_pav2.crc_inst.crc5_q[0] ),
    .B1_N(_08480_),
    .X(_01189_));
 a41o_1 _13093_ (.A1(\digitop_pav2.crc_inst.count[2] ),
    .A2(\digitop_pav2.crc_inst.count[1] ),
    .A3(\digitop_pav2.crc_inst.count[0] ),
    .A4(\digitop_pav2.crc_inst.mctrl_data_end_ff ),
    .B1(\digitop_pav2.crc_inst.count[3] ),
    .X(_01188_));
 nand4_1 _13094_ (.A(\digitop_pav2.crc_inst.count[3] ),
    .B(\digitop_pav2.crc_inst.count[2] ),
    .C(\digitop_pav2.crc_inst.count[1] ),
    .D(\digitop_pav2.crc_inst.count[0] ),
    .Y(_08482_));
 and2_1 _13095_ (.A(\digitop_pav2.crc_inst.mctrl_data_end_ff ),
    .B(_08482_),
    .X(_08483_));
 and3_1 _13096_ (.A(\digitop_pav2.crc_inst.count[1] ),
    .B(\digitop_pav2.crc_inst.count[0] ),
    .C(_08483_),
    .X(_08484_));
 xor2_1 _13097_ (.A(\digitop_pav2.crc_inst.count[2] ),
    .B(_08484_),
    .X(_01187_));
 a21oi_1 _13098_ (.A1(\digitop_pav2.crc_inst.count[0] ),
    .A2(\digitop_pav2.crc_inst.mctrl_data_end_ff ),
    .B1(\digitop_pav2.crc_inst.count[1] ),
    .Y(_08485_));
 nor2_1 _13099_ (.A(_08484_),
    .B(_08485_),
    .Y(_01186_));
 nor2_1 _13100_ (.A(\digitop_pav2.crc_inst.count[0] ),
    .B(\digitop_pav2.crc_inst.mctrl_data_end_ff ),
    .Y(_08486_));
 a21oi_1 _13101_ (.A1(\digitop_pav2.crc_inst.count[0] ),
    .A2(_08483_),
    .B1(_08486_),
    .Y(_01185_));
 and2_1 _13102_ (.A(\digitop_pav2.crc_eval ),
    .B(_08482_),
    .X(_08487_));
 nor2_1 _13103_ (.A(_07259_),
    .B(_07270_),
    .Y(_08488_));
 or3_1 _13104_ (.A(\digitop_pav2.sec_inst.shift_out.st[7] ),
    .B(net701),
    .C(net707),
    .X(_08489_));
 or2_1 _13105_ (.A(\digitop_pav2.sec_inst.shift_out.st[5] ),
    .B(net709),
    .X(_08490_));
 or2_1 _13106_ (.A(_08489_),
    .B(_08490_),
    .X(_08491_));
 nor2_1 _13107_ (.A(\digitop_pav2.sec_inst.shift_out.st[2] ),
    .B(_08491_),
    .Y(_08492_));
 or3_2 _13108_ (.A(\digitop_pav2.sec_inst.shift_out.st[4] ),
    .B(\digitop_pav2.sec_inst.shift_out.st[7] ),
    .C(\digitop_pav2.sec_inst.shift_out.st[0] ),
    .X(_08493_));
 nor2_1 _13109_ (.A(_08490_),
    .B(_08493_),
    .Y(_08494_));
 nor2_1 _13110_ (.A(net704),
    .B(_08494_),
    .Y(_08495_));
 and2_1 _13111_ (.A(\digitop_pav2.sec_inst.shift_out.ctr[1] ),
    .B(\digitop_pav2.sec_inst.shift_out.ctr[0] ),
    .X(_08496_));
 nand2_1 _13112_ (.A(\digitop_pav2.sec_inst.shift_out.ctr[1] ),
    .B(\digitop_pav2.sec_inst.shift_out.ctr[0] ),
    .Y(_08497_));
 nand2_1 _13113_ (.A(net705),
    .B(_08496_),
    .Y(_08498_));
 a21o_1 _13114_ (.A1(net704),
    .A2(_08494_),
    .B1(_08498_),
    .X(_08499_));
 or2_1 _13115_ (.A(_08495_),
    .B(_08499_),
    .X(_08500_));
 or3_1 _13116_ (.A(\digitop_pav2.sec_inst.shift_out.st[2] ),
    .B(net701),
    .C(net707),
    .X(_08501_));
 a21oi_1 _13117_ (.A1(\digitop_pav2.sec_inst.shift_out.j_ctr[6] ),
    .A2(_08490_),
    .B1(_08501_),
    .Y(_08502_));
 o2bb2a_1 _13118_ (.A1_N(\digitop_pav2.sec_inst.en_shifto ),
    .A2_N(_08492_),
    .B1(_08500_),
    .B2(_08502_),
    .X(_08503_));
 and2b_2 _13119_ (.A_N(\digitop_pav2.sec_inst.shift_out.st[4] ),
    .B(_08503_),
    .X(_08504_));
 inv_2 _13120_ (.A(_08504_),
    .Y(_08505_));
 and2_1 _13121_ (.A(net702),
    .B(net701),
    .X(_08506_));
 nor2_1 _13122_ (.A(\digitop_pav2.sec_inst.shift_out.st[2] ),
    .B(\digitop_pav2.sec_inst.shift_out.st[4] ),
    .Y(_08507_));
 or4_1 _13123_ (.A(\digitop_pav2.sec_inst.shift_out.st[2] ),
    .B(\digitop_pav2.sec_inst.shift_out.st[4] ),
    .C(\digitop_pav2.sec_inst.shift_out.st[5] ),
    .D(\digitop_pav2.sec_inst.shift_out.st[7] ),
    .X(_08508_));
 a21o_1 _13124_ (.A1(net709),
    .A2(_08506_),
    .B1(_08508_),
    .X(_08509_));
 and4_1 _13125_ (.A(\digitop_pav2.ack_inst.cnt_ff[0] ),
    .B(net1182),
    .C(\digitop_pav2.ack_inst.cnt_ff[2] ),
    .D(\digitop_pav2.ack_inst.cnt_ff[3] ),
    .X(_08510_));
 and3_1 _13126_ (.A(\digitop_pav2.ack_inst.rcnt_ff[0] ),
    .B(\digitop_pav2.ack_inst.rcnt_ff[1] ),
    .C(_08510_),
    .X(_08511_));
 nor2_2 _13127_ (.A(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[0] ),
    .B(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[1] ),
    .Y(_08512_));
 or3b_1 _13128_ (.A(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[2] ),
    .B(_07118_),
    .C_N(_08512_),
    .X(_08513_));
 inv_2 _13129_ (.A(_08513_),
    .Y(_08514_));
 a221o_1 _13130_ (.A1(\digitop_pav2.ack_inst.g_ack_i ),
    .A2(_08511_),
    .B1(_08514_),
    .B2(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[4] ),
    .C1(\digitop_pav2.access_inst.access_ctrl0.dt_acc_done_o ),
    .X(_08515_));
 a31o_2 _13131_ (.A1(_08491_),
    .A2(_08505_),
    .A3(_08509_),
    .B1(_08515_),
    .X(_08516_));
 and2_1 _13132_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[5] ),
    .B(_08516_),
    .X(_08517_));
 o31a_1 _13133_ (.A1(net1181),
    .A2(_07260_),
    .A3(_07291_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[5] ),
    .X(_08518_));
 a21o_1 _13134_ (.A1(_08516_),
    .A2(_08518_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[12] ),
    .X(_08519_));
 o21a_2 _13135_ (.A1(_08487_),
    .A2(_08519_),
    .B1(\digitop_pav2.crc_inst.dt_tx_en_aux ),
    .X(_08520_));
 or2_1 _13136_ (.A(net1302),
    .B(_08520_),
    .X(_08521_));
 inv_2 _13137_ (.A(net525),
    .Y(_08522_));
 mux2_1 _13138_ (.A0(\digitop_pav2.crc_inst.crc16_q[15] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[14] ),
    .S(net525),
    .X(_01165_));
 mux2_1 _13139_ (.A0(\digitop_pav2.crc_inst.crc16_q[14] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[13] ),
    .S(net525),
    .X(_01164_));
 mux2_1 _13140_ (.A0(\digitop_pav2.crc_inst.crc16_q[13] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[12] ),
    .S(net524),
    .X(_01163_));
 nor2_1 _13141_ (.A(net1296),
    .B(_07071_),
    .Y(_08523_));
 nand2_1 _13142_ (.A(_07121_),
    .B(_08507_),
    .Y(_08524_));
 nor3_1 _13143_ (.A(\digitop_pav2.sec_inst.shift_out.st[5] ),
    .B(_08489_),
    .C(_08524_),
    .Y(_08525_));
 and2_1 _13144_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[4] ),
    .B(net582),
    .X(_08526_));
 nand2_1 _13145_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[4] ),
    .B(net582),
    .Y(_08527_));
 and2_1 _13146_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[3] ),
    .B(net582),
    .X(_08528_));
 nand2_1 _13147_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[3] ),
    .B(net582),
    .Y(_08529_));
 nand2_1 _13148_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[0] ),
    .B(net582),
    .Y(_08530_));
 nand2_1 _13149_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[1] ),
    .B(net582),
    .Y(_08531_));
 mux2_1 _13150_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[105] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[121] ),
    .S(net564),
    .X(_08532_));
 nand2_1 _13151_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[2] ),
    .B(net582),
    .Y(_08533_));
 mux2_1 _13152_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[89] ),
    .A1(_08532_),
    .S(net562),
    .X(_08534_));
 mux2_1 _13153_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[73] ),
    .A1(_08534_),
    .S(net560),
    .X(_08535_));
 mux2_1 _13154_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[57] ),
    .A1(_08535_),
    .S(net566),
    .X(_08536_));
 and2_1 _13155_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[5] ),
    .B(net582),
    .X(_08537_));
 nand2_1 _13156_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[5] ),
    .B(net582),
    .Y(_08538_));
 a21o_1 _13157_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[41] ),
    .A2(_08526_),
    .B1(_08537_),
    .X(_08539_));
 a21o_1 _13158_ (.A1(net568),
    .A2(_08536_),
    .B1(_08539_),
    .X(_08540_));
 and2_1 _13159_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[6] ),
    .B(net582),
    .X(_08541_));
 nand2_1 _13160_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[6] ),
    .B(_08525_),
    .Y(_08542_));
 o21a_1 _13161_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[25] ),
    .A2(net558),
    .B1(net556),
    .X(_08543_));
 a221o_1 _13162_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[9] ),
    .A2(_08541_),
    .B1(_08543_),
    .B2(_08540_),
    .C1(net700),
    .X(_08544_));
 nor3_1 _13163_ (.A(net709),
    .B(_08489_),
    .C(_08524_),
    .Y(_08545_));
 and2_1 _13164_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[4] ),
    .B(net580),
    .X(_08546_));
 nand2_1 _13165_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[4] ),
    .B(net580),
    .Y(_08547_));
 nand2_1 _13166_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[3] ),
    .B(net580),
    .Y(_08548_));
 nor2_1 _13167_ (.A(net366),
    .B(net552),
    .Y(_08549_));
 and2_1 _13168_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[0] ),
    .B(net580),
    .X(_08550_));
 nand2_1 _13169_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[0] ),
    .B(net580),
    .Y(_08551_));
 and2_1 _13170_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[1] ),
    .B(net580),
    .X(_08552_));
 nand2_1 _13171_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[1] ),
    .B(net580),
    .Y(_08553_));
 mux2_1 _13172_ (.A0(_08172_),
    .A1(_08173_),
    .S(net549),
    .X(_08554_));
 and2_1 _13173_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[2] ),
    .B(net580),
    .X(_08555_));
 nand2_1 _13174_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[2] ),
    .B(net580),
    .Y(_08556_));
 nor2_1 _13175_ (.A(net366),
    .B(net544),
    .Y(_08557_));
 a221o_1 _13176_ (.A1(net544),
    .A2(_08554_),
    .B1(_08557_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[9] ),
    .C1(net543),
    .X(_08558_));
 a21o_1 _13177_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[9] ),
    .A2(net370),
    .B1(net541),
    .X(_08559_));
 a32o_1 _13178_ (.A1(net551),
    .A2(_08558_),
    .A3(_08559_),
    .B1(net336),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[9] ),
    .X(_08560_));
 and2_2 _13179_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[5] ),
    .B(net580),
    .X(_08561_));
 nand2_1 _13180_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[5] ),
    .B(net581),
    .Y(_08562_));
 a31o_1 _13181_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[9] ),
    .A2(net372),
    .A3(net555),
    .B1(_08561_),
    .X(_08563_));
 a21o_1 _13182_ (.A1(net553),
    .A2(_08560_),
    .B1(_08563_),
    .X(_08564_));
 and2_2 _13183_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[6] ),
    .B(net581),
    .X(_08565_));
 nand2_1 _13184_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[6] ),
    .B(net581),
    .Y(_08566_));
 a21o_1 _13185_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[9] ),
    .A2(net372),
    .B1(net539),
    .X(_08567_));
 a21o_1 _13186_ (.A1(_08178_),
    .A2(_08565_),
    .B1(net708),
    .X(_08568_));
 a31o_1 _13187_ (.A1(_08564_),
    .A2(net538),
    .A3(_08567_),
    .B1(_08568_),
    .X(_08569_));
 and2b_1 _13188_ (.A_N(net703),
    .B(net705),
    .X(_08570_));
 and2b_2 _13189_ (.A_N(\digitop_pav2.sec_inst.shift_out.ctr[0] ),
    .B(\digitop_pav2.sec_inst.shift_out.ctr[1] ),
    .X(_08571_));
 and4_1 _13190_ (.A(_08544_),
    .B(_08569_),
    .C(_08570_),
    .D(_08571_),
    .X(_08572_));
 mux2_1 _13191_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[97] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[113] ),
    .S(net564),
    .X(_08573_));
 mux2_1 _13192_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[81] ),
    .A1(_08573_),
    .S(net562),
    .X(_08574_));
 mux2_1 _13193_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[65] ),
    .A1(_08574_),
    .S(net560),
    .X(_08575_));
 mux2_1 _13194_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[49] ),
    .A1(_08575_),
    .S(net566),
    .X(_08576_));
 mux2_1 _13195_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[33] ),
    .A1(_08576_),
    .S(net568),
    .X(_08577_));
 mux2_1 _13196_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[17] ),
    .A1(_08577_),
    .S(net558),
    .X(_08578_));
 mux2_1 _13197_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[1] ),
    .A1(_08578_),
    .S(net556),
    .X(_08579_));
 a21o_1 _13198_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[1] ),
    .A2(net379),
    .B1(net547),
    .X(_08580_));
 a21o_1 _13199_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[1] ),
    .A2(net379),
    .B1(net549),
    .X(_08581_));
 a31o_1 _13200_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[1] ),
    .A2(net379),
    .A3(_08552_),
    .B1(net543),
    .X(_08582_));
 a31o_1 _13201_ (.A1(net544),
    .A2(_08580_),
    .A3(_08581_),
    .B1(_08582_),
    .X(_08583_));
 a21o_1 _13202_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[1] ),
    .A2(net379),
    .B1(net541),
    .X(_08584_));
 a32o_1 _13203_ (.A1(net551),
    .A2(_08583_),
    .A3(_08584_),
    .B1(net336),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[1] ),
    .X(_08585_));
 nor2_1 _13204_ (.A(net366),
    .B(net553),
    .Y(_08586_));
 a221o_1 _13205_ (.A1(net554),
    .A2(_08585_),
    .B1(_08586_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[1] ),
    .C1(_08561_),
    .X(_08587_));
 o211a_1 _13206_ (.A1(_08279_),
    .A2(net539),
    .B1(net537),
    .C1(_08587_),
    .X(_08588_));
 a311o_1 _13207_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[1] ),
    .A2(net386),
    .A3(_08565_),
    .B1(_08588_),
    .C1(net709),
    .X(_08589_));
 and3_1 _13208_ (.A(net703),
    .B(net705),
    .C(_08571_),
    .X(_08590_));
 o211a_1 _13209_ (.A1(net699),
    .A2(_08579_),
    .B1(_08589_),
    .C1(_08590_),
    .X(_08591_));
 mux2_1 _13210_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[104] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[120] ),
    .S(net564),
    .X(_08592_));
 mux2_1 _13211_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[88] ),
    .A1(_08592_),
    .S(net562),
    .X(_08593_));
 mux2_1 _13212_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[72] ),
    .A1(_08593_),
    .S(net560),
    .X(_08594_));
 mux2_1 _13213_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[56] ),
    .A1(_08594_),
    .S(net566),
    .X(_08595_));
 mux2_1 _13214_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[40] ),
    .A1(_08595_),
    .S(net568),
    .X(_08596_));
 mux2_1 _13215_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[24] ),
    .A1(_08596_),
    .S(net558),
    .X(_08597_));
 mux2_1 _13216_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[8] ),
    .A1(_08597_),
    .S(net556),
    .X(_08598_));
 a21o_1 _13217_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[8] ),
    .A2(net369),
    .B1(net547),
    .X(_08599_));
 a21o_1 _13218_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[8] ),
    .A2(net369),
    .B1(net549),
    .X(_08600_));
 a31o_1 _13219_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[8] ),
    .A2(net369),
    .A3(net546),
    .B1(net543),
    .X(_08601_));
 a31o_1 _13220_ (.A1(net544),
    .A2(_08599_),
    .A3(_08600_),
    .B1(_08601_),
    .X(_08602_));
 a21o_1 _13221_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[8] ),
    .A2(net369),
    .B1(net541),
    .X(_08603_));
 a32o_1 _13222_ (.A1(net551),
    .A2(_08602_),
    .A3(_08603_),
    .B1(net336),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[8] ),
    .X(_08604_));
 a31o_1 _13223_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[8] ),
    .A2(net372),
    .A3(net555),
    .B1(_08561_),
    .X(_08605_));
 a21o_1 _13224_ (.A1(net553),
    .A2(_08604_),
    .B1(_08605_),
    .X(_08606_));
 a21o_1 _13225_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[8] ),
    .A2(net372),
    .B1(net539),
    .X(_08607_));
 o21ai_1 _13226_ (.A1(_08346_),
    .A2(net538),
    .B1(net700),
    .Y(_08608_));
 a31o_1 _13227_ (.A1(net538),
    .A2(_08606_),
    .A3(_08607_),
    .B1(_08608_),
    .X(_08609_));
 nor2_1 _13228_ (.A(net703),
    .B(_08498_),
    .Y(_08610_));
 o211a_1 _13229_ (.A1(net699),
    .A2(_08598_),
    .B1(_08609_),
    .C1(_08610_),
    .X(_08611_));
 a21o_1 _13230_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[2] ),
    .A2(net378),
    .B1(net549),
    .X(_08612_));
 a21o_1 _13231_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[2] ),
    .A2(net377),
    .B1(net547),
    .X(_08613_));
 a31o_1 _13232_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[2] ),
    .A2(net378),
    .A3(net546),
    .B1(net543),
    .X(_08614_));
 a31o_1 _13233_ (.A1(net545),
    .A2(_08612_),
    .A3(_08613_),
    .B1(_08614_),
    .X(_08615_));
 o211a_1 _13234_ (.A1(_08246_),
    .A2(net542),
    .B1(_08615_),
    .C1(net552),
    .X(_08616_));
 a21oi_1 _13235_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[2] ),
    .A2(net336),
    .B1(_08616_),
    .Y(_08617_));
 nor2_1 _13236_ (.A(net555),
    .B(_08617_),
    .Y(_08618_));
 a211o_1 _13237_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[2] ),
    .A2(_08586_),
    .B1(_08618_),
    .C1(_08561_),
    .X(_08619_));
 a21o_1 _13238_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[2] ),
    .A2(net385),
    .B1(net539),
    .X(_08620_));
 nor2_1 _13239_ (.A(net366),
    .B(net537),
    .Y(_08621_));
 a32o_1 _13240_ (.A1(net537),
    .A2(_08619_),
    .A3(_08620_),
    .B1(_08621_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ),
    .X(_08622_));
 mux2_1 _13241_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[98] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[114] ),
    .S(net565),
    .X(_08623_));
 mux2_1 _13242_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[82] ),
    .A1(_08623_),
    .S(net563),
    .X(_08624_));
 mux2_1 _13243_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[66] ),
    .A1(_08624_),
    .S(net561),
    .X(_08625_));
 mux2_1 _13244_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[50] ),
    .A1(_08625_),
    .S(net567),
    .X(_08626_));
 mux2_1 _13245_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[34] ),
    .A1(_08626_),
    .S(net569),
    .X(_08627_));
 mux2_1 _13246_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[18] ),
    .A1(_08627_),
    .S(net559),
    .X(_08628_));
 mux2_1 _13247_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[2] ),
    .A1(_08628_),
    .S(net557),
    .X(_08629_));
 and2b_2 _13248_ (.A_N(\digitop_pav2.sec_inst.shift_out.ctr[1] ),
    .B(\digitop_pav2.sec_inst.shift_out.ctr[0] ),
    .X(_08630_));
 o2111a_1 _13249_ (.A1(net699),
    .A2(_08629_),
    .B1(_08630_),
    .C1(net704),
    .D1(net705),
    .X(_08631_));
 o21ai_1 _13250_ (.A1(net708),
    .A2(_08622_),
    .B1(_08631_),
    .Y(_08632_));
 nor2_2 _13251_ (.A(\digitop_pav2.sec_inst.shift_out.ctr[1] ),
    .B(\digitop_pav2.sec_inst.shift_out.ctr[0] ),
    .Y(_08633_));
 nor2_1 _13252_ (.A(net704),
    .B(net705),
    .Y(_08634_));
 a21o_1 _13253_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[12] ),
    .A2(net378),
    .B1(net547),
    .X(_08635_));
 a21o_1 _13254_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[12] ),
    .A2(net378),
    .B1(net549),
    .X(_08636_));
 a31o_1 _13255_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[12] ),
    .A2(net381),
    .A3(net546),
    .B1(net543),
    .X(_08637_));
 a31o_1 _13256_ (.A1(net545),
    .A2(_08635_),
    .A3(_08636_),
    .B1(_08637_),
    .X(_08638_));
 a21o_1 _13257_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[12] ),
    .A2(net378),
    .B1(net541),
    .X(_08639_));
 a21o_1 _13258_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[12] ),
    .A2(net336),
    .B1(net555),
    .X(_08640_));
 a31o_1 _13259_ (.A1(net551),
    .A2(_08638_),
    .A3(_08639_),
    .B1(_08640_),
    .X(_08641_));
 a21o_1 _13260_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[12] ),
    .A2(net385),
    .B1(net553),
    .X(_08642_));
 nor2_2 _13261_ (.A(net366),
    .B(net539),
    .Y(_08643_));
 nor2_1 _13262_ (.A(_08298_),
    .B(net538),
    .Y(_08644_));
 a32o_1 _13263_ (.A1(net539),
    .A2(_08641_),
    .A3(_08642_),
    .B1(_08643_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[12] ),
    .X(_08645_));
 a211o_1 _13264_ (.A1(net538),
    .A2(_08645_),
    .B1(_08644_),
    .C1(net708),
    .X(_08646_));
 mux2_1 _13265_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[108] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[124] ),
    .S(net564),
    .X(_08647_));
 mux2_1 _13266_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[92] ),
    .A1(_08647_),
    .S(net562),
    .X(_08648_));
 mux2_1 _13267_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[76] ),
    .A1(_08648_),
    .S(net560),
    .X(_08649_));
 mux2_1 _13268_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[60] ),
    .A1(_08649_),
    .S(net566),
    .X(_08650_));
 mux2_1 _13269_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[44] ),
    .A1(_08650_),
    .S(net568),
    .X(_08651_));
 or2_1 _13270_ (.A(_08537_),
    .B(_08651_),
    .X(_08652_));
 o21a_1 _13271_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[28] ),
    .A2(net558),
    .B1(net556),
    .X(_08653_));
 a221o_1 _13272_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[12] ),
    .A2(_08541_),
    .B1(_08652_),
    .B2(_08653_),
    .C1(net700),
    .X(_08654_));
 nor2_1 _13273_ (.A(net706),
    .B(_08497_),
    .Y(_08655_));
 a21o_1 _13274_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[4] ),
    .A2(net379),
    .B1(net550),
    .X(_08656_));
 a21o_1 _13275_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[4] ),
    .A2(net379),
    .B1(net547),
    .X(_08657_));
 a31o_1 _13276_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[4] ),
    .A2(net379),
    .A3(net546),
    .B1(_08555_),
    .X(_08658_));
 a31o_1 _13277_ (.A1(net545),
    .A2(_08656_),
    .A3(_08657_),
    .B1(_08658_),
    .X(_08659_));
 o211a_1 _13278_ (.A1(_08160_),
    .A2(net542),
    .B1(_08659_),
    .C1(net552),
    .X(_08660_));
 a211o_1 _13279_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[4] ),
    .A2(net337),
    .B1(_08660_),
    .C1(net555),
    .X(_08661_));
 a21o_1 _13280_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[4] ),
    .A2(net385),
    .B1(net554),
    .X(_08662_));
 a32o_1 _13281_ (.A1(net540),
    .A2(_08661_),
    .A3(_08662_),
    .B1(_08643_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[4] ),
    .X(_08663_));
 a221o_1 _13282_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[4] ),
    .A2(_08621_),
    .B1(_08663_),
    .B2(net537),
    .C1(net708),
    .X(_08664_));
 mux2_1 _13283_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[100] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[116] ),
    .S(net565),
    .X(_08665_));
 mux2_1 _13284_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[84] ),
    .A1(_08665_),
    .S(net563),
    .X(_08666_));
 mux2_1 _13285_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[68] ),
    .A1(_08666_),
    .S(net561),
    .X(_08667_));
 mux2_1 _13286_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[52] ),
    .A1(_08667_),
    .S(net567),
    .X(_08668_));
 mux2_1 _13287_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[36] ),
    .A1(_08668_),
    .S(net569),
    .X(_08669_));
 mux2_1 _13288_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[20] ),
    .A1(_08669_),
    .S(net559),
    .X(_08670_));
 mux2_1 _13289_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[4] ),
    .A1(_08670_),
    .S(net557),
    .X(_08671_));
 o2111a_1 _13290_ (.A1(net699),
    .A2(_08671_),
    .B1(_08664_),
    .C1(_08655_),
    .D1(net703),
    .X(_08672_));
 mux2_1 _13291_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[110] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[126] ),
    .S(net564),
    .X(_08673_));
 mux2_1 _13292_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[94] ),
    .A1(_08673_),
    .S(net562),
    .X(_08674_));
 mux2_1 _13293_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[78] ),
    .A1(_08674_),
    .S(net560),
    .X(_08675_));
 or2_1 _13294_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[62] ),
    .B(net566),
    .X(_08676_));
 o211a_1 _13295_ (.A1(_08528_),
    .A2(_08675_),
    .B1(_08676_),
    .C1(net568),
    .X(_08677_));
 a211o_1 _13296_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[46] ),
    .A2(_08526_),
    .B1(_08537_),
    .C1(_08677_),
    .X(_08678_));
 o21a_1 _13297_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[30] ),
    .A2(net558),
    .B1(net556),
    .X(_08679_));
 a221o_1 _13298_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[14] ),
    .A2(_08541_),
    .B1(_08678_),
    .B2(_08679_),
    .C1(net700),
    .X(_08680_));
 a21o_1 _13299_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[14] ),
    .A2(net370),
    .B1(net547),
    .X(_08681_));
 a21o_1 _13300_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[14] ),
    .A2(net370),
    .B1(net549),
    .X(_08682_));
 a31o_1 _13301_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[14] ),
    .A2(net369),
    .A3(net546),
    .B1(net543),
    .X(_08683_));
 a31o_1 _13302_ (.A1(net544),
    .A2(_08681_),
    .A3(_08682_),
    .B1(_08683_),
    .X(_08684_));
 a21o_1 _13303_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[14] ),
    .A2(net369),
    .B1(net541),
    .X(_08685_));
 a21o_1 _13304_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[14] ),
    .A2(net336),
    .B1(net555),
    .X(_08686_));
 a31o_1 _13305_ (.A1(net551),
    .A2(_08684_),
    .A3(_08685_),
    .B1(_08686_),
    .X(_08687_));
 o211a_1 _13306_ (.A1(_08388_),
    .A2(net553),
    .B1(net539),
    .C1(_08687_),
    .X(_08688_));
 a31o_1 _13307_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[14] ),
    .A2(net372),
    .A3(_08561_),
    .B1(_08565_),
    .X(_08689_));
 o22a_1 _13308_ (.A1(_08393_),
    .A2(net538),
    .B1(_08688_),
    .B2(_08689_),
    .X(_08690_));
 o211a_1 _13309_ (.A1(net708),
    .A2(_08690_),
    .B1(_08634_),
    .C1(_08630_),
    .X(_08691_));
 mux2_1 _13310_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[109] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[125] ),
    .S(net564),
    .X(_08692_));
 mux2_1 _13311_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[93] ),
    .A1(_08692_),
    .S(net562),
    .X(_08693_));
 mux2_1 _13312_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[77] ),
    .A1(_08693_),
    .S(net560),
    .X(_08694_));
 mux2_1 _13313_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[61] ),
    .A1(_08694_),
    .S(net566),
    .X(_08695_));
 mux2_1 _13314_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[45] ),
    .A1(_08695_),
    .S(net568),
    .X(_08696_));
 mux2_1 _13315_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[29] ),
    .A1(_08696_),
    .S(net558),
    .X(_08697_));
 mux2_1 _13316_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[13] ),
    .A1(_08697_),
    .S(net556),
    .X(_08698_));
 a21o_1 _13317_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[13] ),
    .A2(net377),
    .B1(net548),
    .X(_08699_));
 a21o_1 _13318_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[13] ),
    .A2(net377),
    .B1(net550),
    .X(_08700_));
 a31o_1 _13319_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[13] ),
    .A2(net377),
    .A3(net546),
    .B1(net543),
    .X(_08701_));
 a31o_1 _13320_ (.A1(net544),
    .A2(_08699_),
    .A3(_08700_),
    .B1(_08701_),
    .X(_08702_));
 a21o_1 _13321_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[13] ),
    .A2(net377),
    .B1(net542),
    .X(_08703_));
 a32o_1 _13322_ (.A1(net552),
    .A2(_08702_),
    .A3(_08703_),
    .B1(net337),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[13] ),
    .X(_08704_));
 a221o_1 _13323_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[13] ),
    .A2(_08586_),
    .B1(_08704_),
    .B2(net553),
    .C1(_08561_),
    .X(_08705_));
 o211a_1 _13324_ (.A1(_08190_),
    .A2(net540),
    .B1(net537),
    .C1(_08705_),
    .X(_08706_));
 a21o_1 _13325_ (.A1(_08196_),
    .A2(_08565_),
    .B1(net708),
    .X(_08707_));
 o22a_1 _13326_ (.A1(net699),
    .A2(_08698_),
    .B1(_08706_),
    .B2(_08707_),
    .X(_08708_));
 nor2_1 _13327_ (.A(net366),
    .B(net541),
    .Y(_08709_));
 a31o_1 _13328_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[0] ),
    .A2(net380),
    .A3(net548),
    .B1(_08552_),
    .X(_08710_));
 a31o_1 _13329_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[0] ),
    .A2(net379),
    .A3(net550),
    .B1(_08710_),
    .X(_08711_));
 a21o_1 _13330_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[0] ),
    .A2(net380),
    .B1(net545),
    .X(_08712_));
 a32o_1 _13331_ (.A1(net542),
    .A2(_08711_),
    .A3(_08712_),
    .B1(_08709_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ),
    .X(_08713_));
 a22o_1 _13332_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[0] ),
    .A2(net337),
    .B1(_08713_),
    .B2(net551),
    .X(_08714_));
 a31o_1 _13333_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[0] ),
    .A2(net386),
    .A3(net555),
    .B1(_08561_),
    .X(_08715_));
 a21o_1 _13334_ (.A1(net554),
    .A2(_08714_),
    .B1(_08715_),
    .X(_08716_));
 o211a_1 _13335_ (.A1(_08311_),
    .A2(net540),
    .B1(net537),
    .C1(_08716_),
    .X(_08717_));
 a31o_1 _13336_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[0] ),
    .A2(net386),
    .A3(_08565_),
    .B1(net709),
    .X(_08718_));
 mux2_1 _13337_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[96] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[112] ),
    .S(net565),
    .X(_08719_));
 mux2_1 _13338_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[80] ),
    .A1(_08719_),
    .S(net563),
    .X(_08720_));
 mux2_1 _13339_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[64] ),
    .A1(_08720_),
    .S(net561),
    .X(_08721_));
 mux2_1 _13340_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[48] ),
    .A1(_08721_),
    .S(net567),
    .X(_08722_));
 mux2_1 _13341_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[32] ),
    .A1(_08722_),
    .S(net569),
    .X(_08723_));
 mux2_1 _13342_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[16] ),
    .A1(_08723_),
    .S(net559),
    .X(_08724_));
 mux2_1 _13343_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[0] ),
    .A1(_08724_),
    .S(net557),
    .X(_08725_));
 o22a_1 _13344_ (.A1(_08717_),
    .A2(_08718_),
    .B1(_08725_),
    .B2(net699),
    .X(_08726_));
 and4_1 _13345_ (.A(net703),
    .B(net705),
    .C(_08496_),
    .D(_08726_),
    .X(_08727_));
 mux2_1 _13346_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[101] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[117] ),
    .S(net565),
    .X(_08728_));
 mux2_1 _13347_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[85] ),
    .A1(_08728_),
    .S(net563),
    .X(_08729_));
 mux2_1 _13348_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[69] ),
    .A1(_08729_),
    .S(net561),
    .X(_08730_));
 mux2_1 _13349_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[53] ),
    .A1(_08730_),
    .S(net567),
    .X(_08731_));
 mux2_1 _13350_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[37] ),
    .A1(_08731_),
    .S(net569),
    .X(_08732_));
 mux2_1 _13351_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[21] ),
    .A1(_08732_),
    .S(net559),
    .X(_08733_));
 and3b_1 _13352_ (.A_N(net705),
    .B(_08571_),
    .C(net703),
    .X(_08734_));
 mux2_1 _13353_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[102] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[118] ),
    .S(net565),
    .X(_08735_));
 mux2_1 _13354_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[86] ),
    .A1(_08735_),
    .S(net563),
    .X(_08736_));
 mux2_1 _13355_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[70] ),
    .A1(_08736_),
    .S(net561),
    .X(_08737_));
 mux2_1 _13356_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[54] ),
    .A1(_08737_),
    .S(net567),
    .X(_08738_));
 mux2_1 _13357_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[38] ),
    .A1(_08738_),
    .S(net569),
    .X(_08739_));
 mux2_1 _13358_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[22] ),
    .A1(_08739_),
    .S(net559),
    .X(_08740_));
 and3b_1 _13359_ (.A_N(net705),
    .B(_08630_),
    .C(net703),
    .X(_08741_));
 a31o_1 _13360_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ),
    .A2(net385),
    .A3(_08565_),
    .B1(net708),
    .X(_08742_));
 and3_1 _13361_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ),
    .B(net377),
    .C(net543),
    .X(_08743_));
 a31o_1 _13362_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[7] ),
    .A2(net377),
    .A3(net549),
    .B1(net546),
    .X(_08744_));
 a31o_1 _13363_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[7] ),
    .A2(net370),
    .A3(net547),
    .B1(_08744_),
    .X(_08745_));
 a21o_1 _13364_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ),
    .A2(net377),
    .B1(net544),
    .X(_08746_));
 a31o_1 _13365_ (.A1(net541),
    .A2(_08745_),
    .A3(_08746_),
    .B1(_08743_),
    .X(_08747_));
 a22o_1 _13366_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[7] ),
    .A2(net336),
    .B1(_08747_),
    .B2(net551),
    .X(_08748_));
 a22o_1 _13367_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[7] ),
    .A2(_08586_),
    .B1(_08748_),
    .B2(net553),
    .X(_08749_));
 a22o_1 _13368_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ),
    .A2(_08643_),
    .B1(_08749_),
    .B2(net539),
    .X(_08750_));
 a21o_1 _13369_ (.A1(net538),
    .A2(_08750_),
    .B1(_08742_),
    .X(_08751_));
 mux2_1 _13370_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[103] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[119] ),
    .S(net564),
    .X(_08752_));
 mux2_1 _13371_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[87] ),
    .A1(_08752_),
    .S(net562),
    .X(_08753_));
 mux2_1 _13372_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[71] ),
    .A1(_08753_),
    .S(net560),
    .X(_08754_));
 or2_1 _13373_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[55] ),
    .B(net566),
    .X(_08755_));
 o211a_1 _13374_ (.A1(_08528_),
    .A2(_08754_),
    .B1(_08755_),
    .C1(net568),
    .X(_08756_));
 a211o_1 _13375_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[39] ),
    .A2(_08526_),
    .B1(_08537_),
    .C1(_08756_),
    .X(_08757_));
 o21a_1 _13376_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[23] ),
    .A2(net558),
    .B1(net556),
    .X(_08758_));
 a221o_1 _13377_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[7] ),
    .A2(_08541_),
    .B1(_08757_),
    .B2(_08758_),
    .C1(net700),
    .X(_08759_));
 and4b_1 _13378_ (.A_N(net705),
    .B(_08633_),
    .C(_08759_),
    .D(net703),
    .X(_08760_));
 mux2_1 _13379_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[99] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[115] ),
    .S(net565),
    .X(_08761_));
 mux2_1 _13380_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[83] ),
    .A1(_08761_),
    .S(net563),
    .X(_08762_));
 mux2_1 _13381_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[67] ),
    .A1(_08762_),
    .S(net561),
    .X(_08763_));
 mux2_1 _13382_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[51] ),
    .A1(_08763_),
    .S(net567),
    .X(_08764_));
 mux2_1 _13383_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[35] ),
    .A1(_08764_),
    .S(net569),
    .X(_08765_));
 mux2_1 _13384_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[19] ),
    .A1(_08765_),
    .S(net559),
    .X(_08766_));
 mux2_1 _13385_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[3] ),
    .A1(_08766_),
    .S(net557),
    .X(_08767_));
 a21o_1 _13386_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[3] ),
    .A2(net377),
    .B1(net542),
    .X(_08768_));
 and3_1 _13387_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[3] ),
    .B(net377),
    .C(net550),
    .X(_08769_));
 a31o_1 _13388_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[3] ),
    .A2(net378),
    .A3(net548),
    .B1(_08769_),
    .X(_08770_));
 a221o_1 _13389_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[3] ),
    .A2(_08557_),
    .B1(_08770_),
    .B2(net545),
    .C1(_08555_),
    .X(_08771_));
 a21o_1 _13390_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[3] ),
    .A2(net337),
    .B1(net555),
    .X(_08772_));
 a31o_1 _13391_ (.A1(net552),
    .A2(_08768_),
    .A3(_08771_),
    .B1(_08772_),
    .X(_08773_));
 a21o_1 _13392_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[3] ),
    .A2(net385),
    .B1(net554),
    .X(_08774_));
 a21o_1 _13393_ (.A1(_08773_),
    .A2(_08774_),
    .B1(_08561_),
    .X(_08775_));
 a21o_1 _13394_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[3] ),
    .A2(net385),
    .B1(net540),
    .X(_08776_));
 o21ai_1 _13395_ (.A1(_08138_),
    .A2(_08566_),
    .B1(net699),
    .Y(_08777_));
 a31o_1 _13396_ (.A1(net537),
    .A2(_08775_),
    .A3(_08776_),
    .B1(_08777_),
    .X(_08778_));
 o2111a_1 _13397_ (.A1(net699),
    .A2(_08767_),
    .B1(_08633_),
    .C1(net706),
    .D1(net703),
    .X(_08779_));
 a21o_1 _13398_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[11] ),
    .A2(net369),
    .B1(net549),
    .X(_08780_));
 a21o_1 _13399_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[11] ),
    .A2(net369),
    .B1(net547),
    .X(_08781_));
 a31o_1 _13400_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[11] ),
    .A2(net369),
    .A3(net546),
    .B1(net543),
    .X(_08782_));
 a31o_1 _13401_ (.A1(net544),
    .A2(_08780_),
    .A3(_08781_),
    .B1(_08782_),
    .X(_08783_));
 a21o_1 _13402_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[11] ),
    .A2(net369),
    .B1(net541),
    .X(_08784_));
 a32o_1 _13403_ (.A1(net551),
    .A2(_08783_),
    .A3(_08784_),
    .B1(net336),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[11] ),
    .X(_08785_));
 a221o_1 _13404_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[11] ),
    .A2(_08586_),
    .B1(_08785_),
    .B2(net553),
    .C1(_08561_),
    .X(_08786_));
 a21o_1 _13405_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[11] ),
    .A2(net372),
    .B1(net539),
    .X(_08787_));
 a21o_1 _13406_ (.A1(_08377_),
    .A2(_08565_),
    .B1(net708),
    .X(_08788_));
 a31o_1 _13407_ (.A1(net538),
    .A2(_08786_),
    .A3(_08787_),
    .B1(_08788_),
    .X(_08789_));
 a21o_1 _13408_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[5] ),
    .A2(net380),
    .B1(net550),
    .X(_08790_));
 a21o_1 _13409_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[5] ),
    .A2(net380),
    .B1(net548),
    .X(_08791_));
 a31o_1 _13410_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[5] ),
    .A2(net380),
    .A3(_08552_),
    .B1(_08555_),
    .X(_08792_));
 a31o_1 _13411_ (.A1(net545),
    .A2(_08790_),
    .A3(_08791_),
    .B1(_08792_),
    .X(_08793_));
 o211a_1 _13412_ (.A1(_08359_),
    .A2(net542),
    .B1(_08793_),
    .C1(net552),
    .X(_08794_));
 a211o_1 _13413_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[5] ),
    .A2(net337),
    .B1(_08794_),
    .C1(_08546_),
    .X(_08795_));
 a21o_1 _13414_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[5] ),
    .A2(net385),
    .B1(net554),
    .X(_08796_));
 and3_1 _13415_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[6] ),
    .B(net379),
    .C(net550),
    .X(_08797_));
 a31o_1 _13416_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[6] ),
    .A2(net379),
    .A3(net548),
    .B1(_08797_),
    .X(_08798_));
 a221o_1 _13417_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[6] ),
    .A2(_08557_),
    .B1(_08798_),
    .B2(net545),
    .C1(_08555_),
    .X(_08799_));
 a21o_1 _13418_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[6] ),
    .A2(net380),
    .B1(net542),
    .X(_08800_));
 a21o_1 _13419_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[6] ),
    .A2(net337),
    .B1(_08546_),
    .X(_08801_));
 a31o_1 _13420_ (.A1(net552),
    .A2(_08799_),
    .A3(_08800_),
    .B1(_08801_),
    .X(_08802_));
 o211a_1 _13421_ (.A1(_08208_),
    .A2(net554),
    .B1(net540),
    .C1(_08802_),
    .X(_08803_));
 a31o_1 _13422_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[10] ),
    .A2(net378),
    .A3(net547),
    .B1(net546),
    .X(_08804_));
 a31o_1 _13423_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ),
    .A2(net378),
    .A3(net549),
    .B1(_08804_),
    .X(_08805_));
 a21o_1 _13424_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[10] ),
    .A2(net378),
    .B1(net544),
    .X(_08806_));
 a32o_1 _13425_ (.A1(net541),
    .A2(_08805_),
    .A3(_08806_),
    .B1(_08709_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ),
    .X(_08807_));
 and2_1 _13426_ (.A(net551),
    .B(_08807_),
    .X(_08808_));
 a211o_1 _13427_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[10] ),
    .A2(net336),
    .B1(_08808_),
    .C1(net555),
    .X(_08809_));
 a21o_1 _13428_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[10] ),
    .A2(net385),
    .B1(net553),
    .X(_08810_));
 a32o_1 _13429_ (.A1(net540),
    .A2(_08809_),
    .A3(_08810_),
    .B1(_08643_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[10] ),
    .X(_08811_));
 nor2_1 _13430_ (.A(_08265_),
    .B(net537),
    .Y(_08812_));
 a211o_1 _13431_ (.A1(net537),
    .A2(_08811_),
    .B1(_08812_),
    .C1(net708),
    .X(_08813_));
 mux2_1 _13432_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[106] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[122] ),
    .S(net564),
    .X(_08814_));
 mux2_1 _13433_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[90] ),
    .A1(_08814_),
    .S(net562),
    .X(_08815_));
 mux2_1 _13434_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[74] ),
    .A1(_08815_),
    .S(net560),
    .X(_08816_));
 mux2_1 _13435_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[58] ),
    .A1(_08816_),
    .S(net566),
    .X(_08817_));
 mux2_1 _13436_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[42] ),
    .A1(_08817_),
    .S(net568),
    .X(_08818_));
 mux2_1 _13437_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[26] ),
    .A1(_08818_),
    .S(net558),
    .X(_08819_));
 mux2_1 _13438_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[10] ),
    .A1(_08819_),
    .S(net556),
    .X(_08820_));
 o2111a_1 _13439_ (.A1(net699),
    .A2(_08820_),
    .B1(_08813_),
    .C1(_08630_),
    .D1(_08570_),
    .X(_08821_));
 mux2_1 _13440_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[107] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[123] ),
    .S(net564),
    .X(_08822_));
 mux2_1 _13441_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[91] ),
    .A1(_08822_),
    .S(net562),
    .X(_08823_));
 mux2_1 _13442_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[75] ),
    .A1(_08823_),
    .S(net560),
    .X(_08824_));
 mux2_1 _13443_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[59] ),
    .A1(_08824_),
    .S(net566),
    .X(_08825_));
 a21o_1 _13444_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[43] ),
    .A2(_08526_),
    .B1(_08537_),
    .X(_08826_));
 a21o_1 _13445_ (.A1(net568),
    .A2(_08825_),
    .B1(_08826_),
    .X(_08827_));
 mux2_1 _13446_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[5] ),
    .A1(_08733_),
    .S(net557),
    .X(_08828_));
 a32o_1 _13447_ (.A1(net540),
    .A2(_08795_),
    .A3(_08796_),
    .B1(_08643_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[5] ),
    .X(_08829_));
 a221o_1 _13448_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[5] ),
    .A2(_08621_),
    .B1(_08829_),
    .B2(net537),
    .C1(net708),
    .X(_08830_));
 o211a_1 _13449_ (.A1(net699),
    .A2(_08828_),
    .B1(_08830_),
    .C1(_08734_),
    .X(_08831_));
 o21a_1 _13450_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[27] ),
    .A2(net558),
    .B1(net556),
    .X(_08832_));
 a221o_1 _13451_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[11] ),
    .A2(_08541_),
    .B1(_08827_),
    .B2(_08832_),
    .C1(net700),
    .X(_08833_));
 and4_1 _13452_ (.A(_08570_),
    .B(_08633_),
    .C(_08789_),
    .D(_08833_),
    .X(_08834_));
 a21oi_1 _13453_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[6] ),
    .A2(_08643_),
    .B1(_08803_),
    .Y(_08835_));
 nor2_1 _13454_ (.A(_08565_),
    .B(_08835_),
    .Y(_08836_));
 a211o_1 _13455_ (.A1(_08213_),
    .A2(_08565_),
    .B1(_08836_),
    .C1(net709),
    .X(_08837_));
 mux2_1 _13456_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[6] ),
    .A1(_08740_),
    .S(net557),
    .X(_08838_));
 o211a_1 _13457_ (.A1(net700),
    .A2(_08838_),
    .B1(_08837_),
    .C1(_08741_),
    .X(_08839_));
 a41o_1 _13458_ (.A1(_08496_),
    .A2(_08634_),
    .A3(_08646_),
    .A4(_08654_),
    .B1(_08821_),
    .X(_08840_));
 or4b_1 _13459_ (.A(_08572_),
    .B(_08591_),
    .C(_08611_),
    .D_N(_08632_),
    .X(_08841_));
 or4_1 _13460_ (.A(_08672_),
    .B(_08834_),
    .C(_08839_),
    .D(_08841_),
    .X(_08842_));
 a221o_1 _13461_ (.A1(_08633_),
    .A2(_08634_),
    .B1(_08778_),
    .B2(_08779_),
    .C1(_08831_),
    .X(_08843_));
 a311o_1 _13462_ (.A1(_08571_),
    .A2(_08634_),
    .A3(_08708_),
    .B1(_08727_),
    .C1(_08843_),
    .X(_08844_));
 a211o_1 _13463_ (.A1(_08680_),
    .A2(_08691_),
    .B1(_08842_),
    .C1(_08844_),
    .X(_08845_));
 a211o_1 _13464_ (.A1(_08751_),
    .A2(_08760_),
    .B1(_08840_),
    .C1(_08845_),
    .X(_08846_));
 nor2_1 _13465_ (.A(net583),
    .B(net581),
    .Y(_08847_));
 mux2_1 _13466_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[111] ),
    .A1(\digitop_pav2.sec_inst.r128.reg128_o[127] ),
    .S(net564),
    .X(_08848_));
 mux2_1 _13467_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[95] ),
    .A1(_08848_),
    .S(net562),
    .X(_08849_));
 mux2_1 _13468_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[79] ),
    .A1(_08849_),
    .S(net560),
    .X(_08850_));
 mux2_1 _13469_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[63] ),
    .A1(_08850_),
    .S(net566),
    .X(_08851_));
 mux2_1 _13470_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[47] ),
    .A1(_08851_),
    .S(net568),
    .X(_08852_));
 mux2_1 _13471_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[31] ),
    .A1(_08852_),
    .S(net558),
    .X(_08853_));
 mux2_1 _13472_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[15] ),
    .A1(_08853_),
    .S(net556),
    .X(_08854_));
 a21o_1 _13473_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[15] ),
    .A2(net370),
    .B1(net547),
    .X(_08855_));
 a21o_1 _13474_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[15] ),
    .A2(net370),
    .B1(net549),
    .X(_08856_));
 a31o_1 _13475_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[15] ),
    .A2(net370),
    .A3(net546),
    .B1(net543),
    .X(_08857_));
 a31o_1 _13476_ (.A1(net544),
    .A2(_08855_),
    .A3(_08856_),
    .B1(_08857_),
    .X(_08858_));
 a21o_1 _13477_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[15] ),
    .A2(net370),
    .B1(net541),
    .X(_08859_));
 a32o_1 _13478_ (.A1(net551),
    .A2(_08858_),
    .A3(_08859_),
    .B1(net336),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[15] ),
    .X(_08860_));
 a31o_1 _13479_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[15] ),
    .A2(net372),
    .A3(net555),
    .B1(_08561_),
    .X(_08861_));
 a21o_1 _13480_ (.A1(net553),
    .A2(_08860_),
    .B1(_08861_),
    .X(_08862_));
 a21o_1 _13481_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[15] ),
    .A2(net372),
    .B1(net539),
    .X(_08863_));
 o21ai_1 _13482_ (.A1(_08234_),
    .A2(net538),
    .B1(net700),
    .Y(_08864_));
 a31o_1 _13483_ (.A1(net538),
    .A2(_08862_),
    .A3(_08863_),
    .B1(_08864_),
    .X(_08865_));
 o21a_1 _13484_ (.A1(net700),
    .A2(_08854_),
    .B1(_08865_),
    .X(_08866_));
 or4b_1 _13485_ (.A(net703),
    .B(net705),
    .C(_08866_),
    .D_N(_08633_),
    .X(_08867_));
 a21o_1 _13486_ (.A1(_08846_),
    .A2(_08867_),
    .B1(_08847_),
    .X(_08868_));
 o311a_1 _13487_ (.A1(net583),
    .A2(net581),
    .A3(_08726_),
    .B1(_08868_),
    .C1(_08490_),
    .X(_08869_));
 nor3_4 _13488_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[6] ),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[5] ),
    .C(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[1] ),
    .Y(_08870_));
 or3_2 _13489_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[6] ),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[5] ),
    .C(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[1] ),
    .X(_08871_));
 nand2_1 _13490_ (.A(net1650),
    .B(_07334_),
    .Y(_08872_));
 nor2_2 _13491_ (.A(_08870_),
    .B(_08872_),
    .Y(_08873_));
 or2_2 _13492_ (.A(_08870_),
    .B(_08872_),
    .X(_08874_));
 nor2_1 _13493_ (.A(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[2] ),
    .B(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[3] ),
    .Y(_08875_));
 a21oi_1 _13494_ (.A1(_08512_),
    .A2(_08875_),
    .B1(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[4] ),
    .Y(_08876_));
 and2_2 _13495_ (.A(net1475),
    .B(net1736),
    .X(_08877_));
 and2b_1 _13496_ (.A_N(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[1] ),
    .B(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[0] ),
    .X(_08878_));
 nand2_1 _13497_ (.A(net1474),
    .B(\digitop_pav2.func_rng_data[15] ),
    .Y(_08879_));
 inv_2 _13498_ (.A(_08879_),
    .Y(_08880_));
 and2_2 _13499_ (.A(net1474),
    .B(net1776),
    .X(_08881_));
 and2b_1 _13500_ (.A_N(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[0] ),
    .B(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[1] ),
    .X(_08882_));
 and2_2 _13501_ (.A(net1476),
    .B(net1781),
    .X(_08883_));
 a22o_1 _13502_ (.A1(_08878_),
    .A2(_08880_),
    .B1(_08882_),
    .B2(_08883_),
    .X(_08884_));
 a31o_1 _13503_ (.A1(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[0] ),
    .A2(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[1] ),
    .A3(_08881_),
    .B1(_08884_),
    .X(_08885_));
 and2_1 _13504_ (.A(net1474),
    .B(\digitop_pav2.func_rng_data[3] ),
    .X(_08886_));
 nand2_1 _13505_ (.A(net1474),
    .B(net1741),
    .Y(_08887_));
 and3_1 _13506_ (.A(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[0] ),
    .B(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[1] ),
    .C(_08886_),
    .X(_08888_));
 and2_2 _13507_ (.A(net1475),
    .B(net1734),
    .X(_08889_));
 and2_2 _13508_ (.A(net1475),
    .B(net1765),
    .X(_08890_));
 and2_2 _13509_ (.A(net1475),
    .B(net1766),
    .X(_08891_));
 a221o_1 _13510_ (.A1(_08512_),
    .A2(_08889_),
    .B1(_08890_),
    .B2(_08882_),
    .C1(_08888_),
    .X(_08892_));
 a21o_1 _13511_ (.A1(_08878_),
    .A2(_08891_),
    .B1(_08892_),
    .X(_08893_));
 and3b_1 _13512_ (.A_N(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[2] ),
    .B(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[3] ),
    .C(_08893_),
    .X(_08894_));
 and2_2 _13513_ (.A(net1770),
    .B(net1474),
    .X(_08895_));
 nand2_1 _13514_ (.A(\digitop_pav2.func_rng_data[5] ),
    .B(net1474),
    .Y(_08896_));
 and2_1 _13515_ (.A(net1476),
    .B(\digitop_pav2.func_rng_data[7] ),
    .X(_08897_));
 nand2_1 _13516_ (.A(net1476),
    .B(\digitop_pav2.func_rng_data[7] ),
    .Y(_08898_));
 a22o_1 _13517_ (.A1(_08882_),
    .A2(_08895_),
    .B1(_08897_),
    .B2(_08878_),
    .X(_08899_));
 and2_2 _13518_ (.A(net1476),
    .B(net1768),
    .X(_08900_));
 nand2_1 _13519_ (.A(net1476),
    .B(\digitop_pav2.func_rng_data[6] ),
    .Y(_08901_));
 and3_1 _13520_ (.A(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[0] ),
    .B(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[1] ),
    .C(_08900_),
    .X(_08902_));
 and2_2 _13521_ (.A(net1475),
    .B(net1782),
    .X(_08903_));
 nand2_1 _13522_ (.A(net1474),
    .B(\digitop_pav2.func_rng_data[8] ),
    .Y(_08904_));
 a211o_1 _13523_ (.A1(_08512_),
    .A2(_08903_),
    .B1(_08902_),
    .C1(_08899_),
    .X(_08905_));
 a31o_1 _13524_ (.A1(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[2] ),
    .A2(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[3] ),
    .A3(_08905_),
    .B1(_08894_),
    .X(_08906_));
 a21o_1 _13525_ (.A1(_08875_),
    .A2(_08885_),
    .B1(_08906_),
    .X(_08907_));
 and2_2 _13526_ (.A(net1475),
    .B(net1767),
    .X(_08908_));
 and2_2 _13527_ (.A(net1474),
    .B(net1769),
    .X(_08909_));
 a22o_1 _13528_ (.A1(_08878_),
    .A2(_08908_),
    .B1(_08909_),
    .B2(_08882_),
    .X(_08910_));
 and2_2 _13529_ (.A(net1474),
    .B(net1780),
    .X(_08911_));
 nand2_1 _13530_ (.A(net1474),
    .B(\digitop_pav2.func_rng_data[9] ),
    .Y(_08912_));
 and2_2 _13531_ (.A(net1475),
    .B(net1806),
    .X(_08913_));
 and3_1 _13532_ (.A(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[0] ),
    .B(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[1] ),
    .C(_08913_),
    .X(_08914_));
 a211o_1 _13533_ (.A1(_08512_),
    .A2(_08911_),
    .B1(_08914_),
    .C1(_08910_),
    .X(_08915_));
 a31o_1 _13534_ (.A1(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[2] ),
    .A2(_07118_),
    .A3(_08915_),
    .B1(_08907_),
    .X(_08916_));
 mux2_1 _13535_ (.A0(_08877_),
    .A1(_08916_),
    .S(_08876_),
    .X(_08917_));
 a31o_1 _13536_ (.A1(\digitop_pav2.ack_inst.cnt_ff[0] ),
    .A2(net1182),
    .A3(\digitop_pav2.ack_inst.buffer_ff[8] ),
    .B1(\digitop_pav2.ack_inst.cnt_ff[3] ),
    .X(_08918_));
 nor2_1 _13537_ (.A(_07054_),
    .B(net1182),
    .Y(_08919_));
 and2_1 _13538_ (.A(_07054_),
    .B(net1182),
    .X(_08920_));
 nor2_1 _13539_ (.A(\digitop_pav2.ack_inst.cnt_ff[0] ),
    .B(net1182),
    .Y(_08921_));
 a221o_1 _13540_ (.A1(\digitop_pav2.ack_inst.buffer_ff[9] ),
    .A2(_08920_),
    .B1(_08921_),
    .B2(\digitop_pav2.ack_inst.buffer_ff[11] ),
    .C1(_08918_),
    .X(_08922_));
 a21o_1 _13541_ (.A1(\digitop_pav2.ack_inst.buffer_ff[10] ),
    .A2(_08919_),
    .B1(_08922_),
    .X(_08923_));
 and3_1 _13542_ (.A(\digitop_pav2.ack_inst.cnt_ff[0] ),
    .B(net1182),
    .C(\digitop_pav2.ack_inst.buffer_ff[0] ),
    .X(_08924_));
 a221o_1 _13543_ (.A1(\digitop_pav2.ack_inst.buffer_ff[2] ),
    .A2(_08919_),
    .B1(_08920_),
    .B2(\digitop_pav2.ack_inst.buffer_ff[1] ),
    .C1(_08924_),
    .X(_08925_));
 a211o_1 _13544_ (.A1(\digitop_pav2.ack_inst.buffer_ff[3] ),
    .A2(_08921_),
    .B1(_08925_),
    .C1(_07089_),
    .X(_08926_));
 a2111o_1 _13545_ (.A1(_07036_),
    .A2(\digitop_pav2.access_inst.access_ctrl0.state[15] ),
    .B1(net1142),
    .C1(net1143),
    .D1(\digitop_pav2.access_inst.access_ctrl0.state[22] ),
    .X(_08927_));
 a32o_1 _13546_ (.A1(_07121_),
    .A2(\digitop_pav2.fg_tc ),
    .A3(_08492_),
    .B1(_08927_),
    .B2(\digitop_pav2.access_inst.access_ctrl0.tx_bit_i ),
    .X(_08928_));
 and3_1 _13547_ (.A(\digitop_pav2.ack_inst.cnt_ff[0] ),
    .B(\digitop_pav2.ack_inst.cnt_ff[1] ),
    .C(\digitop_pav2.ack_inst.buffer_ff[12] ),
    .X(_08929_));
 a221o_1 _13548_ (.A1(_07054_),
    .A2(\digitop_pav2.ack_inst.buffer_ff[13] ),
    .B1(\digitop_pav2.ack_inst.buffer_ff[14] ),
    .B2(_08919_),
    .C1(_08921_),
    .X(_08930_));
 o32a_1 _13549_ (.A1(\digitop_pav2.ack_inst.cnt_ff[0] ),
    .A2(net1182),
    .A3(\digitop_pav2.ack_inst.buffer_ff[15] ),
    .B1(_08929_),
    .B2(_08930_),
    .X(_08931_));
 and3_1 _13550_ (.A(\digitop_pav2.ack_inst.cnt_ff[0] ),
    .B(net1182),
    .C(\digitop_pav2.ack_inst.buffer_ff[4] ),
    .X(_08932_));
 a221o_1 _13551_ (.A1(\digitop_pav2.ack_inst.buffer_ff[6] ),
    .A2(_08919_),
    .B1(_08921_),
    .B2(\digitop_pav2.ack_inst.buffer_ff[7] ),
    .C1(_08932_),
    .X(_08933_));
 a211o_1 _13552_ (.A1(\digitop_pav2.ack_inst.buffer_ff[5] ),
    .A2(_08920_),
    .B1(_08933_),
    .C1(_07089_),
    .X(_08934_));
 o211a_1 _13553_ (.A1(\digitop_pav2.ack_inst.cnt_ff[3] ),
    .A2(_08931_),
    .B1(_08934_),
    .C1(_07088_),
    .X(_08935_));
 a31o_1 _13554_ (.A1(\digitop_pav2.ack_inst.cnt_ff[2] ),
    .A2(_08923_),
    .A3(_08926_),
    .B1(_08928_),
    .X(_08936_));
 a22o_1 _13555_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[13] ),
    .A2(_08571_),
    .B1(_08630_),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[14] ),
    .X(_08937_));
 or2_1 _13556_ (.A(net706),
    .B(_08633_),
    .X(_08938_));
 a22o_1 _13557_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[5] ),
    .A2(_08571_),
    .B1(_08630_),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[6] ),
    .X(_08939_));
 a221o_1 _13558_ (.A1(net707),
    .A2(_08937_),
    .B1(_08939_),
    .B2(net701),
    .C1(_08938_),
    .X(_08940_));
 a22o_1 _13559_ (.A1(net701),
    .A2(\digitop_pav2.access_inst.access_transceiver0.handle_i[3] ),
    .B1(\digitop_pav2.access_inst.access_transceiver0.handle_i[11] ),
    .B2(net707),
    .X(_08941_));
 a22o_1 _13560_ (.A1(net701),
    .A2(\digitop_pav2.access_inst.access_transceiver0.handle_i[1] ),
    .B1(\digitop_pav2.access_inst.access_transceiver0.handle_i[9] ),
    .B2(net707),
    .X(_08942_));
 o21ai_1 _13561_ (.A1(net701),
    .A2(net707),
    .B1(net706),
    .Y(_08943_));
 a221o_1 _13562_ (.A1(_08633_),
    .A2(_08941_),
    .B1(_08942_),
    .B2(_08571_),
    .C1(_08943_),
    .X(_08944_));
 a22o_1 _13563_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[8] ),
    .A2(_08496_),
    .B1(_08630_),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[10] ),
    .X(_08945_));
 a22o_1 _13564_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[0] ),
    .A2(_08496_),
    .B1(_08630_),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[2] ),
    .X(_08946_));
 a22o_1 _13565_ (.A1(net707),
    .A2(_08945_),
    .B1(_08946_),
    .B2(net701),
    .X(_08947_));
 o21a_1 _13566_ (.A1(_08944_),
    .A2(_08947_),
    .B1(_08940_),
    .X(_08948_));
 a22o_1 _13567_ (.A1(\digitop_pav2.sec_inst.shift_out.st[1] ),
    .A2(\digitop_pav2.access_inst.access_transceiver0.handle_i[4] ),
    .B1(\digitop_pav2.access_inst.access_transceiver0.handle_i[12] ),
    .B2(net707),
    .X(_08949_));
 a21bo_1 _13568_ (.A1(_08655_),
    .A2(_08949_),
    .B1_N(_08494_),
    .X(_08950_));
 o31a_1 _13569_ (.A1(\digitop_pav2.sec_inst.shift_out.ctr[1] ),
    .A2(\digitop_pav2.sec_inst.shift_out.ctr[0] ),
    .A3(net706),
    .B1(_08494_),
    .X(_08951_));
 a221o_1 _13570_ (.A1(\digitop_pav2.sec_inst.shift_out.st[1] ),
    .A2(\digitop_pav2.access_inst.access_transceiver0.handle_i[7] ),
    .B1(\digitop_pav2.access_inst.access_transceiver0.handle_i[15] ),
    .B2(\digitop_pav2.sec_inst.shift_out.st[6] ),
    .C1(_08951_),
    .X(_08952_));
 o211a_1 _13571_ (.A1(_08948_),
    .A2(_08950_),
    .B1(_08952_),
    .C1(_08501_),
    .X(_08953_));
 a211o_1 _13572_ (.A1(_08873_),
    .A2(_08917_),
    .B1(_08953_),
    .C1(_08869_),
    .X(_08954_));
 or3_2 _13573_ (.A(_08935_),
    .B(_08936_),
    .C(_08954_),
    .X(_08955_));
 a31o_1 _13574_ (.A1(net1296),
    .A2(_08520_),
    .A3(_08955_),
    .B1(_08523_),
    .X(_08956_));
 xnor2_1 _13575_ (.A(_07043_),
    .B(_08956_),
    .Y(_08957_));
 and3b_1 _13576_ (.A_N(_08483_),
    .B(net525),
    .C(_08957_),
    .X(_08958_));
 mux2_1 _13577_ (.A0(\digitop_pav2.crc_inst.crc16_q[12] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[11] ),
    .S(net524),
    .X(_08959_));
 mux2_1 _13578_ (.A0(_08959_),
    .A1(_07044_),
    .S(_08958_),
    .X(_01162_));
 mux2_1 _13579_ (.A0(\digitop_pav2.crc_inst.crc16_q[11] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[10] ),
    .S(net524),
    .X(_01161_));
 mux2_1 _13580_ (.A0(\digitop_pav2.crc_inst.crc16_q[10] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[9] ),
    .S(net524),
    .X(_01160_));
 mux2_1 _13581_ (.A0(\digitop_pav2.crc_inst.crc16_q[9] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[8] ),
    .S(net524),
    .X(_01159_));
 mux2_1 _13582_ (.A0(\digitop_pav2.crc_inst.crc16_q[8] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[7] ),
    .S(net524),
    .X(_01158_));
 mux2_1 _13583_ (.A0(\digitop_pav2.crc_inst.crc16_q[7] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[6] ),
    .S(net525),
    .X(_01157_));
 mux2_1 _13584_ (.A0(\digitop_pav2.crc_inst.crc16_q[6] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[5] ),
    .S(net525),
    .X(_01156_));
 mux2_1 _13585_ (.A0(\digitop_pav2.crc_inst.crc16_q[5] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[4] ),
    .S(net524),
    .X(_08960_));
 mux2_1 _13586_ (.A0(_08960_),
    .A1(_07045_),
    .S(_08958_),
    .X(_01155_));
 mux2_1 _13587_ (.A0(\digitop_pav2.crc_inst.crc16_q[4] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[3] ),
    .S(net525),
    .X(_01154_));
 mux2_1 _13588_ (.A0(\digitop_pav2.crc_inst.crc16_q[3] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[2] ),
    .S(net524),
    .X(_01153_));
 mux2_1 _13589_ (.A0(\digitop_pav2.crc_inst.crc16_q[2] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[1] ),
    .S(net524),
    .X(_01152_));
 mux2_1 _13590_ (.A0(\digitop_pav2.crc_inst.crc16_q[1] ),
    .A1(\digitop_pav2.crc_inst.crc16_q[0] ),
    .S(net524),
    .X(_01151_));
 a21o_1 _13591_ (.A1(\digitop_pav2.crc_inst.crc16_q[0] ),
    .A2(_08522_),
    .B1(_08958_),
    .X(_01150_));
 or2_1 _13592_ (.A(net1453),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_i ),
    .X(_00265_));
 nand2_1 _13593_ (.A(net1399),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_i ),
    .Y(_00264_));
 o211a_1 _13594_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[3] ),
    .A2(_07129_),
    .B1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[4] ),
    .C1(net1273),
    .X(_08961_));
 or3_1 _13595_ (.A(_07063_),
    .B(_07128_),
    .C(_07129_),
    .X(_08962_));
 mux2_1 _13596_ (.A0(_08962_),
    .A1(\digitop_pav2.invent_inst.invent_sel_pav2.mask_mismatch_ff ),
    .S(_08961_),
    .X(_08963_));
 o211a_1 _13597_ (.A1(net1179),
    .A2(net1180),
    .B1(\digitop_pav2.dr ),
    .C1(net1272),
    .X(_08964_));
 and3b_1 _13598_ (.A_N(_08964_),
    .B(_08963_),
    .C(\digitop_pav2.invent_inst.invent_sel_pav2.state[10] ),
    .X(_08965_));
 nor2_1 _13599_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.flags_en_o ),
    .B(net974),
    .Y(_08966_));
 or2_2 _13600_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.flags_en_o ),
    .B(net974),
    .X(_08967_));
 mux2_1 _13601_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[1] ),
    .A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[6] ),
    .S(net1274),
    .X(_08968_));
 mux2_1 _13602_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[0] ),
    .A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[7] ),
    .S(net1274),
    .X(_08969_));
 and2b_1 _13603_ (.A_N(_08969_),
    .B(_08968_),
    .X(_08970_));
 mux2_1 _13604_ (.A0(_07047_),
    .A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_i ),
    .S(_08970_),
    .X(_08971_));
 or2_1 _13605_ (.A(net974),
    .B(_08971_),
    .X(_08972_));
 and2_2 _13606_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[3] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[4] ),
    .X(_08973_));
 and3_1 _13607_ (.A(net1272),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[5] ),
    .C(_08973_),
    .X(_08974_));
 nand2b_2 _13608_ (.A_N(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[4] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[3] ),
    .Y(_08975_));
 or3b_1 _13609_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[3] ),
    .B(_07129_),
    .C_N(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[4] ),
    .X(_08976_));
 a211o_1 _13610_ (.A1(_08975_),
    .A2(_08976_),
    .B1(_07063_),
    .C1(\digitop_pav2.invent_inst.invent_sel_pav2.mask_mismatch_ff ),
    .X(_08977_));
 a31o_1 _13611_ (.A1(net1272),
    .A2(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[3] ),
    .A3(_07129_),
    .B1(_07128_),
    .X(_08978_));
 o31a_1 _13612_ (.A1(_07063_),
    .A2(\digitop_pav2.invent_inst.invent_sel_pav2.mask_mismatch_ff ),
    .A3(_08975_),
    .B1(_08978_),
    .X(_08979_));
 nor2_1 _13613_ (.A(_08974_),
    .B(_08979_),
    .Y(_08980_));
 and3b_1 _13614_ (.A_N(net1179),
    .B(net1180),
    .C(net1272),
    .X(_08981_));
 nand2_1 _13615_ (.A(_08977_),
    .B(_08978_),
    .Y(_08982_));
 inv_2 _13616_ (.A(_08982_),
    .Y(_08983_));
 o21ba_1 _13617_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_i ),
    .A2(_08983_),
    .B1_N(_08980_),
    .X(_08984_));
 o21ai_1 _13618_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_i ),
    .A2(_08981_),
    .B1(net974),
    .Y(_08985_));
 a21o_1 _13619_ (.A1(_08981_),
    .A2(_08984_),
    .B1(_08985_),
    .X(_08986_));
 a21oi_1 _13620_ (.A1(_08972_),
    .A2(_08986_),
    .B1(_08966_),
    .Y(_08987_));
 o21ba_1 _13621_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_r_ff_i ),
    .A2(_08967_),
    .B1_N(_08987_),
    .X(_01092_));
 nand2_1 _13622_ (.A(net1398),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ),
    .Y(_00262_));
 or2_1 _13623_ (.A(net1453),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ),
    .X(_00261_));
 nand2_1 _13624_ (.A(_08968_),
    .B(_08969_),
    .Y(_08988_));
 mux2_1 _13625_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ),
    .A1(_07046_),
    .S(_08988_),
    .X(_08989_));
 a21oi_1 _13626_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.flags_en_o ),
    .A2(_08989_),
    .B1(net975),
    .Y(_08990_));
 a31o_1 _13627_ (.A1(net1272),
    .A2(net1179),
    .A3(net1180),
    .B1(_08964_),
    .X(_08991_));
 o21ai_1 _13628_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ),
    .A2(_08983_),
    .B1(_08991_),
    .Y(_08992_));
 o221a_1 _13629_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ),
    .A2(_08991_),
    .B1(_08992_),
    .B2(_08980_),
    .C1(net975),
    .X(_08993_));
 nor2_1 _13630_ (.A(_08990_),
    .B(_08993_),
    .Y(_08994_));
 a21oi_1 _13631_ (.A1(_07046_),
    .A2(_08966_),
    .B1(_08994_),
    .Y(_01091_));
 a21o_1 _13632_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_s_ff_i ),
    .A2(_08966_),
    .B1(_08987_),
    .X(_01089_));
 or2_1 _13633_ (.A(net1451),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.sl_i ),
    .X(_00256_));
 nand2_1 _13634_ (.A(net1398),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.sl_i ),
    .Y(_00255_));
 or4b_1 _13635_ (.A(_07063_),
    .B(net1179),
    .C(net1180),
    .D_N(\digitop_pav2.dr ),
    .X(_08995_));
 a21oi_1 _13636_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.sl_i ),
    .A2(_08982_),
    .B1(_08980_),
    .Y(_08996_));
 mux2_1 _13637_ (.A0(_08996_),
    .A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.sl_i ),
    .S(_08995_),
    .X(_08997_));
 nor2_1 _13638_ (.A(\digitop_pav2.invent_inst.sl_r_ff ),
    .B(net975),
    .Y(_08998_));
 a21oi_1 _13639_ (.A1(net975),
    .A2(_08997_),
    .B1(_08998_),
    .Y(_01088_));
 mux2_1 _13640_ (.A0(\digitop_pav2.invent_inst.sl_s_ff ),
    .A1(_08997_),
    .S(net975),
    .X(_01087_));
 a21o_1 _13641_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_r_ff_i ),
    .A2(_08966_),
    .B1(_08994_),
    .X(_01078_));
 nand2_1 _13642_ (.A(net1398),
    .B(\digitop_pav2.invent_inst.s1_i ),
    .Y(_00247_));
 or2_1 _13643_ (.A(net1452),
    .B(\digitop_pav2.invent_inst.s1_i ),
    .X(_00246_));
 and3_1 _13644_ (.A(net1274),
    .B(net1247),
    .C(net818),
    .X(_08999_));
 a211o_1 _13645_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[0] ),
    .A2(_08999_),
    .B1(_08967_),
    .C1(\digitop_pav2.invent_inst.invent_sel_pav2.select_valid_o ),
    .X(_09000_));
 and2b_1 _13646_ (.A_N(_08968_),
    .B(_08969_),
    .X(_09001_));
 o21a_1 _13647_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s1_i ),
    .A2(_08977_),
    .B1(_08979_),
    .X(_09002_));
 or4bb_1 _13648_ (.A(_07063_),
    .B(net1180),
    .C_N(net974),
    .D_N(net1179),
    .X(_09003_));
 nand2_1 _13649_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.mask_mismatch_ff ),
    .B(_08974_),
    .Y(_09004_));
 a311o_1 _13650_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s1_i ),
    .A2(\digitop_pav2.invent_inst.invent_sel_pav2.mask_mismatch_ff ),
    .A3(_08974_),
    .B1(_09002_),
    .C1(_09003_),
    .X(_09005_));
 nand2_1 _13651_ (.A(_08967_),
    .B(_09005_),
    .Y(_09006_));
 a21bo_1 _13652_ (.A1(\digitop_pav2.invent_inst.s1_i ),
    .A2(_08966_),
    .B1_N(_09005_),
    .X(_09007_));
 a31o_1 _13653_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.flags_en_o ),
    .A2(_00170_),
    .A3(_09001_),
    .B1(_09007_),
    .X(_09008_));
 mux2_1 _13654_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.s1_i ),
    .A1(_09008_),
    .S(_09000_),
    .X(_01077_));
 and4_1 _13655_ (.A(net1304),
    .B(_07048_),
    .C(net1291),
    .D(net1217),
    .X(_09009_));
 or2_1 _13656_ (.A(net1251),
    .B(_07299_),
    .X(_09010_));
 nor2_1 _13657_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.cmdctr_end3 ),
    .B(_07299_),
    .Y(_09011_));
 o211a_1 _13658_ (.A1(_07295_),
    .A2(_07360_),
    .B1(_07364_),
    .C1(net1294),
    .X(_09012_));
 nor2_1 _13659_ (.A(_07294_),
    .B(_07352_),
    .Y(_09013_));
 or4_1 _13660_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[7] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[6] ),
    .C(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[5] ),
    .D(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[4] ),
    .X(_09014_));
 nor3_1 _13661_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[3] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[2] ),
    .C(_09014_),
    .Y(_09015_));
 and3b_1 _13662_ (.A_N(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[0] ),
    .B(_09015_),
    .C(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[1] ),
    .X(_09016_));
 nand2_1 _13663_ (.A(net1185),
    .B(net1229),
    .Y(_09017_));
 nor2_1 _13664_ (.A(net1189),
    .B(_09017_),
    .Y(_09018_));
 nor2_1 _13665_ (.A(net1216),
    .B(_07352_),
    .Y(_09019_));
 nor2_1 _13666_ (.A(_07354_),
    .B(_09019_),
    .Y(_09020_));
 inv_2 _13667_ (.A(_09020_),
    .Y(_09021_));
 nor4_1 _13668_ (.A(_09012_),
    .B(_09013_),
    .C(_09018_),
    .D(_09021_),
    .Y(_09022_));
 inv_2 _13669_ (.A(net1015),
    .Y(_09023_));
 and2_2 _13670_ (.A(net1302),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[9] ),
    .X(_09024_));
 nand2_1 _13671_ (.A(net1303),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[9] ),
    .Y(_09025_));
 or3b_2 _13672_ (.A(_07257_),
    .B(net1188),
    .C_N(_07347_),
    .X(_09026_));
 inv_2 _13673_ (.A(_09026_),
    .Y(_09027_));
 and4_1 _13674_ (.A(_09010_),
    .B(net1015),
    .C(_09025_),
    .D(_09026_),
    .X(_09028_));
 a21o_1 _13675_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.par4_en_ff ),
    .A2(_09028_),
    .B1(_09011_),
    .X(_00998_));
 a21o_1 _13676_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.par3_en_ff ),
    .A2(_09028_),
    .B1(_09024_),
    .X(_00974_));
 a21o_1 _13677_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.par2_en_ff ),
    .A2(_09028_),
    .B1(_09027_),
    .X(_00973_));
 a41o_1 _13678_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.par1_en_ff ),
    .A2(_09010_),
    .A3(_09025_),
    .A4(_09026_),
    .B1(_09023_),
    .X(_00972_));
 a22o_1 _13679_ (.A1(_09011_),
    .A2(net1188),
    .B1(_09028_),
    .B2(net1251),
    .X(_00971_));
 and3_1 _13680_ (.A(_07067_),
    .B(_07285_),
    .C(_07287_),
    .X(_09029_));
 nor3_1 _13681_ (.A(net1219),
    .B(_07263_),
    .C(net1230),
    .Y(_09030_));
 or3_2 _13682_ (.A(_07245_),
    .B(_07263_),
    .C(net1230),
    .X(_09031_));
 or2_2 _13683_ (.A(_09029_),
    .B(net1187),
    .X(_09032_));
 or4_4 _13684_ (.A(_07243_),
    .B(net1185),
    .C(_07310_),
    .D(_09032_),
    .X(_09033_));
 inv_2 _13685_ (.A(_09033_),
    .Y(_09034_));
 nor2_1 _13686_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.par3_en_ff ),
    .B(_09025_),
    .Y(_09035_));
 or2_2 _13687_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.par3_en_ff ),
    .B(_09025_),
    .X(_09036_));
 or2_1 _13688_ (.A(net1197),
    .B(_09036_),
    .X(_09037_));
 or4_1 _13689_ (.A(_07259_),
    .B(_07361_),
    .C(_09033_),
    .D(_09036_),
    .X(_09038_));
 o21a_2 _13690_ (.A1(_07301_),
    .A2(_09038_),
    .B1(net1304),
    .X(_09039_));
 nand2b_2 _13691_ (.A_N(_09028_),
    .B(_09039_),
    .Y(_09040_));
 nor2_1 _13692_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.par1_en_ff ),
    .B(net1015),
    .Y(_09041_));
 inv_2 _13693_ (.A(_09041_),
    .Y(_09042_));
 nor2_1 _13694_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.par2_en_ff ),
    .B(_09026_),
    .Y(_09043_));
 or2_1 _13695_ (.A(_09041_),
    .B(_09043_),
    .X(_09044_));
 a21oi_1 _13696_ (.A1(net1197),
    .A2(_09035_),
    .B1(_09044_),
    .Y(_09045_));
 inv_2 _13697_ (.A(_09045_),
    .Y(_09046_));
 nor2_2 _13698_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.par4_en_ff ),
    .B(_09010_),
    .Y(_09047_));
 or3_1 _13699_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[2] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[1] ),
    .C(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[0] ),
    .X(_09048_));
 or2_1 _13700_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[3] ),
    .B(_09048_),
    .X(_09049_));
 or3_1 _13701_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[5] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[4] ),
    .C(_09049_),
    .X(_09050_));
 nor2_1 _13702_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[6] ),
    .B(_09050_),
    .Y(_09051_));
 xnor2_1 _13703_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[7] ),
    .B(_09051_),
    .Y(_09052_));
 nor2_1 _13704_ (.A(_09047_),
    .B(_09052_),
    .Y(_09053_));
 o21a_1 _13705_ (.A1(_09035_),
    .A2(_09053_),
    .B1(_09045_),
    .X(_09054_));
 o22a_1 _13706_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[7] ),
    .A2(_09039_),
    .B1(_09040_),
    .B2(_09054_),
    .X(_00970_));
 a31o_1 _13707_ (.A1(net1252),
    .A2(_07268_),
    .A3(_09041_),
    .B1(_09040_),
    .X(_09055_));
 and2_1 _13708_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[6] ),
    .B(_09050_),
    .X(_09056_));
 nor2_1 _13709_ (.A(_09051_),
    .B(_09056_),
    .Y(_09057_));
 o31a_1 _13710_ (.A1(_09035_),
    .A2(_09047_),
    .A3(_09057_),
    .B1(_09037_),
    .X(_09058_));
 nor2_1 _13711_ (.A(_09044_),
    .B(_09058_),
    .Y(_09059_));
 o22a_1 _13712_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[6] ),
    .A2(_09039_),
    .B1(_09055_),
    .B2(_09059_),
    .X(_00969_));
 o21ai_1 _13713_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[4] ),
    .A2(_09049_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[5] ),
    .Y(_09060_));
 a211o_1 _13714_ (.A1(_09050_),
    .A2(_09060_),
    .B1(_09035_),
    .C1(_09047_),
    .X(_09061_));
 a21oi_1 _13715_ (.A1(_09037_),
    .A2(_09061_),
    .B1(_09044_),
    .Y(_09062_));
 o22a_1 _13716_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[5] ),
    .A2(_09039_),
    .B1(_09055_),
    .B2(_09062_),
    .X(_00968_));
 xnor2_1 _13717_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[4] ),
    .B(_09049_),
    .Y(_09063_));
 nand2_1 _13718_ (.A(net1218),
    .B(_09047_),
    .Y(_09064_));
 o211a_1 _13719_ (.A1(_09047_),
    .A2(_09063_),
    .B1(_09064_),
    .C1(_09036_),
    .X(_09065_));
 nor2_1 _13720_ (.A(_09043_),
    .B(_09065_),
    .Y(_09066_));
 a221o_1 _13721_ (.A1(\digitop_pav2.proc_ctrl_inst.cmd.state[2] ),
    .A2(_09043_),
    .B1(_09066_),
    .B2(_09037_),
    .C1(_09041_),
    .X(_09067_));
 o21ai_1 _13722_ (.A1(_07240_),
    .A2(_09042_),
    .B1(_09067_),
    .Y(_09068_));
 o22a_1 _13723_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[4] ),
    .A2(_09039_),
    .B1(_09040_),
    .B2(_09068_),
    .X(_00967_));
 nand2_1 _13724_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[3] ),
    .B(_09048_),
    .Y(_09069_));
 a21oi_1 _13725_ (.A1(_09049_),
    .A2(_09069_),
    .B1(_09047_),
    .Y(_09070_));
 or3_1 _13726_ (.A(_09035_),
    .B(_09043_),
    .C(_09070_),
    .X(_09071_));
 or3_1 _13727_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.par2_en_ff ),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state[2] ),
    .C(_09026_),
    .X(_09072_));
 or4_1 _13728_ (.A(_07258_),
    .B(net1197),
    .C(net1196),
    .D(_07313_),
    .X(_09073_));
 nor2_1 _13729_ (.A(_09042_),
    .B(_09073_),
    .Y(_09074_));
 a31o_1 _13730_ (.A1(_09042_),
    .A2(_09071_),
    .A3(_09072_),
    .B1(_09074_),
    .X(_09075_));
 o22a_1 _13731_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[3] ),
    .A2(_09039_),
    .B1(_09040_),
    .B2(_09075_),
    .X(_00966_));
 a21oi_1 _13732_ (.A1(_07360_),
    .A2(_09041_),
    .B1(_09040_),
    .Y(_09076_));
 o21ai_1 _13733_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[1] ),
    .A2(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[0] ),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[2] ),
    .Y(_09077_));
 a21o_1 _13734_ (.A1(_09048_),
    .A2(_09077_),
    .B1(_09047_),
    .X(_09078_));
 a31o_1 _13735_ (.A1(_09036_),
    .A2(_09064_),
    .A3(_09078_),
    .B1(_09046_),
    .X(_09079_));
 o2bb2a_1 _13736_ (.A1_N(_09076_),
    .A2_N(_09079_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[2] ),
    .B2(_09039_),
    .X(_00965_));
 xor2_1 _13737_ (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[1] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[0] ),
    .X(_09080_));
 o31a_1 _13738_ (.A1(_09035_),
    .A2(_09047_),
    .A3(_09080_),
    .B1(_09037_),
    .X(_09081_));
 or4_1 _13739_ (.A(_07270_),
    .B(net1185),
    .C(_07361_),
    .D(_09042_),
    .X(_09082_));
 o21ai_1 _13740_ (.A1(_09044_),
    .A2(_09081_),
    .B1(_09082_),
    .Y(_09083_));
 o22a_1 _13741_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[1] ),
    .A2(_09039_),
    .B1(_09040_),
    .B2(_09083_),
    .X(_00964_));
 o211a_1 _13742_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[0] ),
    .A2(_09047_),
    .B1(_09064_),
    .C1(_09036_),
    .X(_09084_));
 o21ai_1 _13743_ (.A1(_09046_),
    .A2(_09084_),
    .B1(_09076_),
    .Y(_09085_));
 o21a_1 _13744_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[0] ),
    .A2(_09039_),
    .B1(_09085_),
    .X(_00963_));
 and2_1 _13745_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[1] ),
    .B(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[0] ),
    .X(_09086_));
 and4bb_2 _13746_ (.A_N(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[3] ),
    .B_N(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[2] ),
    .C(_09086_),
    .D(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[4] ),
    .X(_09087_));
 or2_1 _13747_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.pass_t2_flag ),
    .B(_09087_),
    .X(_00956_));
 and3_1 _13748_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[3] ),
    .B(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[2] ),
    .C(_09086_),
    .X(_09088_));
 nor2_1 _13749_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.piex_dt_rx_en_i ),
    .B(_09088_),
    .Y(_09089_));
 or3_1 _13750_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[4] ),
    .B(\digitop_pav2.proc_ctrl_inst.timeout.ctr.piex_dt_rx_en_i ),
    .C(_09088_),
    .X(_00954_));
 a31o_1 _13751_ (.A1(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[2] ),
    .A2(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[1] ),
    .A3(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[0] ),
    .B1(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[3] ),
    .X(_09090_));
 and2_1 _13752_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[4] ),
    .B(_09088_),
    .X(_09091_));
 a221o_1 _13753_ (.A1(\digitop_pav2.proc_ctrl_inst.timeout.ctr.piex_dt_rx_en_i ),
    .A2(_09087_),
    .B1(_09089_),
    .B2(_09090_),
    .C1(_09091_),
    .X(_00953_));
 or2_1 _13754_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[2] ),
    .B(_09086_),
    .X(_09092_));
 a21oi_1 _13755_ (.A1(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[2] ),
    .A2(_09086_),
    .B1(\digitop_pav2.proc_ctrl_inst.timeout.ctr.piex_dt_rx_en_i ),
    .Y(_09093_));
 a221o_1 _13756_ (.A1(\digitop_pav2.proc_ctrl_inst.timeout.ctr.piex_dt_rx_en_i ),
    .A2(_09087_),
    .B1(_09092_),
    .B2(_09093_),
    .C1(_09091_),
    .X(_00952_));
 nor2_1 _13757_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[1] ),
    .B(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[0] ),
    .Y(_09094_));
 nor2_1 _13758_ (.A(_09086_),
    .B(_09094_),
    .Y(_09095_));
 or3_1 _13759_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.piex_dt_rx_en_i ),
    .B(_09091_),
    .C(_09095_),
    .X(_00951_));
 or3b_1 _13760_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.piex_dt_rx_en_i ),
    .B(_09091_),
    .C_N(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[0] ),
    .X(_00950_));
 nor2_1 _13761_ (.A(net1399),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.fm0x_mod_en_i ),
    .Y(_00215_));
 and2b_4 _13762_ (.A_N(net1713),
    .B(net1722),
    .X(_09096_));
 nand2b_4 _13763_ (.A_N(net1713),
    .B(net1722),
    .Y(_09097_));
 a22o_1 _13764_ (.A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[1] ),
    .A2(_08877_),
    .B1(_08881_),
    .B2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[8] ),
    .X(_09098_));
 a221o_1 _13765_ (.A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[5] ),
    .A2(_08886_),
    .B1(_08900_),
    .B2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[11] ),
    .C1(_09098_),
    .X(_09099_));
 a22o_1 _13766_ (.A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[9] ),
    .A2(_08889_),
    .B1(_08909_),
    .B2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[4] ),
    .X(_09100_));
 a221o_1 _13767_ (.A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[3] ),
    .A2(_08897_),
    .B1(_08913_),
    .B2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[6] ),
    .C1(_09100_),
    .X(_09101_));
 a22o_1 _13768_ (.A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[12] ),
    .A2(_08883_),
    .B1(_08891_),
    .B2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[13] ),
    .X(_09102_));
 a221o_1 _13769_ (.A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[15] ),
    .A2(_08895_),
    .B1(_08908_),
    .B2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[14] ),
    .C1(_09102_),
    .X(_09103_));
 a2111o_1 _13770_ (.A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[10] ),
    .A2(_08911_),
    .B1(_09096_),
    .C1(_09101_),
    .D1(_09103_),
    .X(_09104_));
 a22o_1 _13771_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[9] ),
    .A2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[10] ),
    .B1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[12] ),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[13] ),
    .X(_09105_));
 a22o_1 _13772_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[6] ),
    .A2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[11] ),
    .B1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[6] ),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[11] ),
    .X(_09106_));
 a22o_1 _13773_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[3] ),
    .A2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[5] ),
    .B1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[14] ),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[10] ),
    .X(_09107_));
 a221o_1 _13774_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[1] ),
    .A2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[9] ),
    .B1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[15] ),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[5] ),
    .C1(_09107_),
    .X(_09108_));
 a211o_1 _13775_ (.A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[1] ),
    .A2(\digitop_pav2.access_inst.access_transceiver0.handle_i[0] ),
    .B1(_09097_),
    .C1(_09108_),
    .X(_09109_));
 a221o_1 _13776_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[2] ),
    .A2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[13] ),
    .B1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[4] ),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[12] ),
    .C1(_09105_),
    .X(_09110_));
 a221o_1 _13777_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[7] ),
    .A2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[3] ),
    .B1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[8] ),
    .B2(\digitop_pav2.access_inst.access_transceiver0.handle_i[14] ),
    .C1(_09106_),
    .X(_09111_));
 or3_1 _13778_ (.A(_09109_),
    .B(_09110_),
    .C(_09111_),
    .X(_09112_));
 o21a_1 _13779_ (.A1(_09099_),
    .A2(_09104_),
    .B1(_09112_),
    .X(_09113_));
 mux2_1 _13780_ (.A0(\digitop_pav2.access_inst.access_transceiver0.handle_i[4] ),
    .A1(_08890_),
    .S(_09097_),
    .X(_09114_));
 mux2_1 _13781_ (.A0(\digitop_pav2.access_inst.access_transceiver0.handle_i[8] ),
    .A1(_08903_),
    .S(_09097_),
    .X(_09115_));
 or4_1 _13782_ (.A(\digitop_pav2.proc_ctrl_inst.inst_checker.state[15] ),
    .B(\digitop_pav2.proc_ctrl_inst.inst_checker.state[7] ),
    .C(\digitop_pav2.proc_ctrl_inst.inst_checker.state[3] ),
    .D(\digitop_pav2.proc_ctrl_inst.inst_checker.state[11] ),
    .X(_09116_));
 or4_1 _13783_ (.A(\digitop_pav2.proc_ctrl_inst.inst_checker.state[1] ),
    .B(\digitop_pav2.proc_ctrl_inst.inst_checker.state[9] ),
    .C(\digitop_pav2.proc_ctrl_inst.inst_checker.state[5] ),
    .D(\digitop_pav2.proc_ctrl_inst.inst_checker.state[13] ),
    .X(_09117_));
 or4_1 _13784_ (.A(\digitop_pav2.proc_ctrl_inst.inst_checker.state[10] ),
    .B(\digitop_pav2.proc_ctrl_inst.inst_checker.state[2] ),
    .C(\digitop_pav2.proc_ctrl_inst.inst_checker.state[6] ),
    .D(\digitop_pav2.proc_ctrl_inst.inst_checker.state[14] ),
    .X(_09118_));
 or4_1 _13785_ (.A(\digitop_pav2.proc_ctrl_inst.inst_checker.state[12] ),
    .B(\digitop_pav2.proc_ctrl_inst.inst_checker.state[4] ),
    .C(\digitop_pav2.proc_ctrl_inst.inst_checker.state[8] ),
    .D(_09118_),
    .X(_09119_));
 or3_1 _13786_ (.A(_09116_),
    .B(_09117_),
    .C(_09119_),
    .X(_09120_));
 a22o_1 _13787_ (.A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[7] ),
    .A2(_09114_),
    .B1(_09115_),
    .B2(\digitop_pav2.proc_ctrl_inst.inst_checker.state[2] ),
    .X(_09121_));
 or3b_1 _13788_ (.A(_09113_),
    .B(_09121_),
    .C_N(_09120_),
    .X(_09122_));
 mux2_1 _13789_ (.A0(\digitop_pav2.access_inst.access_transceiver0.handle_i[15] ),
    .A1(_08880_),
    .S(_09097_),
    .X(_09123_));
 o21a_1 _13790_ (.A1(_09120_),
    .A2(_09123_),
    .B1(_09122_),
    .X(_09124_));
 xnor2_1 _13791_ (.A(_07071_),
    .B(_09124_),
    .Y(_09125_));
 a21oi_2 _13792_ (.A1(net1167),
    .A2(_09125_),
    .B1(\digitop_pav2.proc_ctrl_inst.inst_checker.dif ),
    .Y(_09126_));
 inv_2 _13793_ (.A(_09126_),
    .Y(_01023_));
 nor2_1 _13794_ (.A(_07274_),
    .B(_01023_),
    .Y(_09127_));
 and4b_1 _13795_ (.A_N(net1249),
    .B(net1293),
    .C(net1186),
    .D(_09127_),
    .X(_09128_));
 or3_1 _13796_ (.A(\digitop_pav2.crc_inst.crc5_q[4] ),
    .B(\digitop_pav2.crc_inst.crc5_q[3] ),
    .C(\digitop_pav2.crc_inst.crc5_q[1] ),
    .X(_09129_));
 or3_1 _13797_ (.A(\digitop_pav2.crc_inst.crc5_q[2] ),
    .B(\digitop_pav2.crc_inst.crc5_q[0] ),
    .C(_09129_),
    .X(_09130_));
 nor2_1 _13798_ (.A(_07048_),
    .B(_09130_),
    .Y(_09131_));
 nand3_1 _13799_ (.A(net1291),
    .B(net1217),
    .C(_09131_),
    .Y(_09132_));
 and4b_1 _13800_ (.A_N(\digitop_pav2.crc_inst.crc16_q[9] ),
    .B(\digitop_pav2.crc_inst.crc16_q[8] ),
    .C(\digitop_pav2.crc_inst.crc16_q[11] ),
    .D(\digitop_pav2.crc_inst.crc16_q[10] ),
    .X(_09133_));
 nor2_1 _13801_ (.A(\digitop_pav2.crc_inst.crc16_q[14] ),
    .B(\digitop_pav2.crc_inst.crc16_q[13] ),
    .Y(_09134_));
 and4_1 _13802_ (.A(_07043_),
    .B(\digitop_pav2.crc_inst.crc16_q[12] ),
    .C(_09133_),
    .D(_09134_),
    .X(_09135_));
 nor4_1 _13803_ (.A(\digitop_pav2.crc_inst.crc16_q[7] ),
    .B(\digitop_pav2.crc_inst.crc16_q[6] ),
    .C(\digitop_pav2.crc_inst.crc16_q[5] ),
    .D(\digitop_pav2.crc_inst.crc16_q[4] ),
    .Y(_09136_));
 and4_1 _13804_ (.A(\digitop_pav2.crc_inst.crc16_q[3] ),
    .B(\digitop_pav2.crc_inst.crc16_q[2] ),
    .C(\digitop_pav2.crc_inst.crc16_q[1] ),
    .D(\digitop_pav2.crc_inst.crc16_q[0] ),
    .X(_09137_));
 nand4_2 _13805_ (.A(net1251),
    .B(_09135_),
    .C(_09136_),
    .D(_09137_),
    .Y(_09138_));
 o41a_1 _13806_ (.A1(net1217),
    .A2(_07297_),
    .A3(net1183),
    .A4(_09138_),
    .B1(_09132_),
    .X(_09139_));
 inv_2 _13807_ (.A(_09139_),
    .Y(_09140_));
 and3_1 _13808_ (.A(net1185),
    .B(_07351_),
    .C(net1189),
    .X(_09141_));
 and2b_1 _13809_ (.A_N(\digitop_pav2.proc_ctrl_inst.cmdfsm.fm0x_dt_tx_st_i ),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[8] ),
    .X(_09142_));
 nor2_2 _13810_ (.A(\digitop_pav2.access_inst.access_ctrl0.replay_nok ),
    .B(\digitop_pav2.access_inst.access_ctrl0.replay_ok ),
    .Y(_09143_));
 or3_2 _13811_ (.A(\digitop_pav2.ack_inst.nvm_ack_rd_stb_o ),
    .B(\digitop_pav2.ack_inst.state_ff[1] ),
    .C(\digitop_pav2.ack_inst.state_ff[2] ),
    .X(_09144_));
 or4_2 _13812_ (.A(\digitop_pav2.access_inst.access_ctrl0.replay_nok ),
    .B(\digitop_pav2.access_inst.access_ctrl0.replay_ok ),
    .C(\digitop_pav2.sec_inst.sm.st[9] ),
    .D(\digitop_pav2.sec_inst.en_shifto ),
    .X(_09145_));
 or3_4 _13813_ (.A(_08871_),
    .B(_09144_),
    .C(_09145_),
    .X(_09146_));
 nor2_1 _13814_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.r_invent3_o ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.r_invent3_o ),
    .Y(_09147_));
 or2_1 _13815_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.r_invent3_o ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.r_invent3_o ),
    .X(_09148_));
 nor2_4 _13816_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.r_invent2_o ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.r_invent2_o ),
    .Y(_09149_));
 nor4_1 _13817_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.r_invent3_o ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.r_invent3_o ),
    .C(\digitop_pav2.invent_inst.invent_qqqr_pav2.r_invent2_o ),
    .D(\digitop_pav2.invent_inst.invent_sel_pav2.r_invent2_o ),
    .Y(_09150_));
 nand2_2 _13818_ (.A(_09147_),
    .B(_09149_),
    .Y(_09151_));
 nor2_1 _13819_ (.A(_09146_),
    .B(_09150_),
    .Y(_09152_));
 or4_4 _13820_ (.A(_08871_),
    .B(_09144_),
    .C(_09145_),
    .D(net1163),
    .X(_09153_));
 o221a_1 _13821_ (.A1(net1217),
    .A2(_07315_),
    .B1(_07332_),
    .B2(_09153_),
    .C1(net1286),
    .X(_09154_));
 or4_1 _13822_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[1] ),
    .B(_09141_),
    .C(_09142_),
    .D(_09154_),
    .X(_09155_));
 nor2_1 _13823_ (.A(\digitop_pav2.crc_inst.crc16_q[6] ),
    .B(\digitop_pav2.crc_inst.crc16_q[5] ),
    .Y(_09156_));
 nor2_1 _13824_ (.A(\digitop_pav2.crc_inst.crc16_q[7] ),
    .B(\digitop_pav2.crc_inst.crc16_q[4] ),
    .Y(_09157_));
 and4_1 _13825_ (.A(_09135_),
    .B(_09137_),
    .C(_09156_),
    .D(_09157_),
    .X(_09158_));
 or3_2 _13826_ (.A(_09128_),
    .B(_09140_),
    .C(_09155_),
    .X(_09159_));
 nand2_1 _13827_ (.A(net1240),
    .B(_07851_),
    .Y(_09160_));
 a31o_1 _13828_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.pass_t1_i ),
    .A2(_09159_),
    .A3(_09160_),
    .B1(\digitop_pav2.sync_inst.inst_clkx.inst_cipher.inst_en.cipher_off_ff ),
    .X(_00582_));
 or4_1 _13829_ (.A(net1051),
    .B(net1053),
    .C(_07600_),
    .D(_07690_),
    .X(_09161_));
 and3b_1 _13830_ (.A_N(net202),
    .B(_07559_),
    .C(_09161_),
    .X(_09162_));
 or4_1 _13831_ (.A(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_crc_en ),
    .B(\digitop_pav2.boot_inst.boot_ctrl0.state[0] ),
    .C(\digitop_pav2.boot_inst.boot_ctrl0.prev_busy ),
    .D(\digitop_pav2.boot_inst.boot_ctrl0.state[3] ),
    .X(_09163_));
 and2_1 _13832_ (.A(net1238),
    .B(net1016),
    .X(_09164_));
 nor2_1 _13833_ (.A(net715),
    .B(net714),
    .Y(_09165_));
 or2_2 _13834_ (.A(net715),
    .B(net714),
    .X(_09166_));
 or4_2 _13835_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[6] ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.state[12] ),
    .C(\digitop_pav2.invent_inst.invent_sel_pav2.state[4] ),
    .D(\digitop_pav2.invent_inst.invent_sel_pav2.state[5] ),
    .X(_09167_));
 a211o_1 _13836_ (.A1(\digitop_pav2.sec_inst.ld_mem.st[0] ),
    .A2(_09166_),
    .B1(_09167_),
    .C1(_09164_),
    .X(_09168_));
 or4b_1 _13837_ (.A(\digitop_pav2.ack_inst.nvm_ack_rd_stb_o ),
    .B(_09162_),
    .C(_09168_),
    .D_N(_09163_),
    .X(_09169_));
 a21o_1 _13838_ (.A1(_07049_),
    .A2(_09169_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.nvm_busy_i ),
    .X(_00577_));
 or3_1 _13839_ (.A(_07283_),
    .B(net1229),
    .C(_07363_),
    .X(_09170_));
 nor4_1 _13840_ (.A(net1290),
    .B(net1295),
    .C(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[6] ),
    .D(net1287),
    .Y(_09171_));
 a22o_1 _13841_ (.A1(_07328_),
    .A2(_09153_),
    .B1(_09170_),
    .B2(net1217),
    .X(_09172_));
 o31a_1 _13842_ (.A1(_07283_),
    .A2(net1229),
    .A3(_07363_),
    .B1(net1215),
    .X(_09173_));
 a21oi_1 _13843_ (.A1(net1217),
    .A2(_09153_),
    .B1(_07087_),
    .Y(_09174_));
 or3b_1 _13844_ (.A(net1304),
    .B(net1251),
    .C_N(net1291),
    .X(_09175_));
 inv_2 _13845_ (.A(_09175_),
    .Y(_09176_));
 a221o_1 _13846_ (.A1(net1296),
    .A2(net1290),
    .B1(net1295),
    .B2(net1183),
    .C1(_09176_),
    .X(_09177_));
 or3_1 _13847_ (.A(_09173_),
    .B(_09174_),
    .C(_09177_),
    .X(_09178_));
 or4_4 _13848_ (.A(net1228),
    .B(_09173_),
    .C(_09174_),
    .D(_09177_),
    .X(_09179_));
 a22oi_4 _13849_ (.A1(\digitop_pav2.pie_inst.fsm.trcal[4] ),
    .A2(net578),
    .B1(net536),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[4] ),
    .Y(_09180_));
 a22oi_1 _13850_ (.A1(\digitop_pav2.memctrl_inst.extra_dt_i[15] ),
    .A2(net578),
    .B1(_09179_),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[3] ),
    .Y(_09181_));
 a22o_1 _13851_ (.A1(\digitop_pav2.memctrl_inst.extra_dt_i[15] ),
    .A2(net579),
    .B1(_09179_),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[3] ),
    .X(_09182_));
 nand2b_1 _13852_ (.A_N(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[2] ),
    .B(net1227),
    .Y(_09183_));
 a221o_1 _13853_ (.A1(\digitop_pav2.memctrl_inst.extra_dt_i[14] ),
    .A2(net578),
    .B1(_09178_),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[2] ),
    .C1(net1227),
    .X(_09184_));
 and3_1 _13854_ (.A(_09182_),
    .B(_09183_),
    .C(_09184_),
    .X(_09185_));
 nand2b_1 _13855_ (.A_N(_09185_),
    .B(_09180_),
    .Y(_09186_));
 a22oi_4 _13856_ (.A1(\digitop_pav2.dr ),
    .A2(net578),
    .B1(net536),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_dr ),
    .Y(_09187_));
 a22o_2 _13857_ (.A1(\digitop_pav2.dr ),
    .A2(net578),
    .B1(net536),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_dr ),
    .X(_09188_));
 nand2b_1 _13858_ (.A_N(_09180_),
    .B(_09185_),
    .Y(_09189_));
 and3_1 _13859_ (.A(_09186_),
    .B(net533),
    .C(_09189_),
    .X(_09190_));
 a22oi_4 _13860_ (.A1(\digitop_pav2.pie_inst.fsm.trcal[6] ),
    .A2(net578),
    .B1(net536),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[6] ),
    .Y(_09191_));
 a22oi_4 _13861_ (.A1(\digitop_pav2.pie_inst.fsm.trcal[7] ),
    .A2(net579),
    .B1(net536),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[7] ),
    .Y(_09192_));
 or2_1 _13862_ (.A(_09191_),
    .B(_09192_),
    .X(_09193_));
 nand2_1 _13863_ (.A(_09191_),
    .B(_09192_),
    .Y(_09194_));
 and2_1 _13864_ (.A(_09193_),
    .B(_09194_),
    .X(_09195_));
 a22oi_4 _13865_ (.A1(\digitop_pav2.pie_inst.fsm.trcal[5] ),
    .A2(net579),
    .B1(net536),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[5] ),
    .Y(_09196_));
 nand2_1 _13866_ (.A(_09191_),
    .B(_09196_),
    .Y(_09197_));
 nor2_1 _13867_ (.A(_09191_),
    .B(_09196_),
    .Y(_09198_));
 or2_1 _13868_ (.A(_09191_),
    .B(_09196_),
    .X(_09199_));
 nor2_1 _13869_ (.A(_09180_),
    .B(_09196_),
    .Y(_09200_));
 or2_1 _13870_ (.A(_09180_),
    .B(_09196_),
    .X(_09201_));
 nand2_1 _13871_ (.A(_09180_),
    .B(_09196_),
    .Y(_09202_));
 nand2_1 _13872_ (.A(_09201_),
    .B(_09202_),
    .Y(_09203_));
 a21oi_1 _13873_ (.A1(_09183_),
    .A2(_09184_),
    .B1(_09182_),
    .Y(_09204_));
 and2_1 _13874_ (.A(_09180_),
    .B(_09181_),
    .X(_09205_));
 o21a_1 _13875_ (.A1(_09173_),
    .A2(_09177_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[0] ),
    .X(_09206_));
 a21o_1 _13876_ (.A1(net1217),
    .A2(_09153_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[0] ),
    .X(_09207_));
 o311a_1 _13877_ (.A1(\digitop_pav2.memctrl_inst.extra_dt_i[12] ),
    .A2(net1215),
    .A3(_09152_),
    .B1(_09207_),
    .C1(net1286),
    .X(_09208_));
 a311o_1 _13878_ (.A1(\digitop_pav2.memctrl_inst.extra_dt_i[12] ),
    .A2(net1217),
    .A3(_09170_),
    .B1(_09206_),
    .C1(_09208_),
    .X(_09209_));
 a22o_1 _13879_ (.A1(\digitop_pav2.memctrl_inst.extra_dt_i[13] ),
    .A2(net578),
    .B1(net536),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[1] ),
    .X(_09210_));
 o221a_1 _13880_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[0] ),
    .A2(_09183_),
    .B1(_09184_),
    .B2(_09209_),
    .C1(_09210_),
    .X(_09211_));
 or4b_2 _13881_ (.A(_09185_),
    .B(_09204_),
    .C(_09205_),
    .D_N(_09211_),
    .X(_09212_));
 o21ba_1 _13882_ (.A1(_09180_),
    .A2(_09181_),
    .B1_N(_09185_),
    .X(_09213_));
 a21o_1 _13883_ (.A1(_09212_),
    .A2(_09213_),
    .B1(_09203_),
    .X(_09214_));
 nand2_2 _13884_ (.A(_09197_),
    .B(_09199_),
    .Y(_09215_));
 a211oi_4 _13885_ (.A1(_09212_),
    .A2(_09213_),
    .B1(_09215_),
    .C1(_09203_),
    .Y(_09216_));
 o31ai_4 _13886_ (.A1(_09198_),
    .A2(_09200_),
    .A3(_09216_),
    .B1(_09195_),
    .Y(_09217_));
 or4_2 _13887_ (.A(_09195_),
    .B(_09198_),
    .C(_09200_),
    .D(_09216_),
    .X(_09218_));
 nand3_1 _13888_ (.A(_09203_),
    .B(_09212_),
    .C(_09213_),
    .Y(_09219_));
 and2_1 _13889_ (.A(_09214_),
    .B(_09219_),
    .X(_09220_));
 and3b_1 _13890_ (.A_N(_09215_),
    .B(_09214_),
    .C(_09201_),
    .X(_09221_));
 a21boi_1 _13891_ (.A1(_09201_),
    .A2(_09214_),
    .B1_N(_09215_),
    .Y(_09222_));
 nand3_1 _13892_ (.A(_09201_),
    .B(_09214_),
    .C(_09215_),
    .Y(_09223_));
 a21o_1 _13893_ (.A1(_09201_),
    .A2(_09214_),
    .B1(_09215_),
    .X(_09224_));
 and3_1 _13894_ (.A(_09220_),
    .B(_09223_),
    .C(_09224_),
    .X(_09225_));
 a32o_1 _13895_ (.A1(_09220_),
    .A2(_09223_),
    .A3(_09224_),
    .B1(_09218_),
    .B2(_09217_),
    .X(_09226_));
 o2111ai_4 _13896_ (.A1(_09221_),
    .A2(_09222_),
    .B1(_09217_),
    .C1(_09218_),
    .D1(_09220_),
    .Y(_09227_));
 a31oi_1 _13897_ (.A1(_09188_),
    .A2(_09226_),
    .A3(_09227_),
    .B1(_09190_),
    .Y(_09228_));
 a31o_2 _13898_ (.A1(_09188_),
    .A2(_09226_),
    .A3(_09227_),
    .B1(_09190_),
    .X(_09229_));
 a22oi_4 _13899_ (.A1(\digitop_pav2.pie_inst.fsm.trcal[8] ),
    .A2(net579),
    .B1(_09179_),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[8] ),
    .Y(_09230_));
 or2_1 _13900_ (.A(_09189_),
    .B(_09199_),
    .X(_09231_));
 or2_1 _13901_ (.A(_09192_),
    .B(_09231_),
    .X(_09232_));
 or2_1 _13902_ (.A(_09192_),
    .B(_09230_),
    .X(_09233_));
 or2_1 _13903_ (.A(_09231_),
    .B(_09233_),
    .X(_09234_));
 nand2_1 _13904_ (.A(_09230_),
    .B(_09232_),
    .Y(_09235_));
 a21o_1 _13905_ (.A1(_09234_),
    .A2(_09235_),
    .B1(_09188_),
    .X(_09236_));
 a22oi_4 _13906_ (.A1(\digitop_pav2.pie_inst.fsm.trcal[9] ),
    .A2(net579),
    .B1(_09179_),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[9] ),
    .Y(_09237_));
 nand2_1 _13907_ (.A(_09192_),
    .B(_09230_),
    .Y(_09238_));
 nand2_1 _13908_ (.A(_09233_),
    .B(_09238_),
    .Y(_09239_));
 inv_2 _13909_ (.A(_09239_),
    .Y(_09240_));
 o311ai_2 _13910_ (.A1(_09198_),
    .A2(_09200_),
    .A3(_09216_),
    .B1(_09240_),
    .C1(_09195_),
    .Y(_09241_));
 and3_1 _13911_ (.A(_09193_),
    .B(_09233_),
    .C(_09241_),
    .X(_09242_));
 a21oi_2 _13912_ (.A1(_09230_),
    .A2(_09242_),
    .B1(_09237_),
    .Y(_09243_));
 and3_1 _13913_ (.A(_09193_),
    .B(_09217_),
    .C(_09239_),
    .X(_09244_));
 a21oi_1 _13914_ (.A1(_09193_),
    .A2(_09217_),
    .B1(_09239_),
    .Y(_09245_));
 or3_2 _13915_ (.A(_09227_),
    .B(_09244_),
    .C(_09245_),
    .X(_09246_));
 nand3b_1 _13916_ (.A_N(_09237_),
    .B(_09242_),
    .C(_09230_),
    .Y(_09247_));
 nor2_2 _13917_ (.A(_09246_),
    .B(_09247_),
    .Y(_09248_));
 o31a_1 _13918_ (.A1(net533),
    .A2(_09243_),
    .A3(_09248_),
    .B1(_09236_),
    .X(_09249_));
 o31ai_4 _13919_ (.A1(net533),
    .A2(_09243_),
    .A3(_09248_),
    .B1(_09236_),
    .Y(_09250_));
 o21ai_1 _13920_ (.A1(_09189_),
    .A2(_09196_),
    .B1(_09191_),
    .Y(_09251_));
 and3_1 _13921_ (.A(net533),
    .B(_09231_),
    .C(_09251_),
    .X(_09252_));
 xor2_1 _13922_ (.A(_09230_),
    .B(_09237_),
    .X(_09253_));
 nand4_1 _13923_ (.A(_09193_),
    .B(_09233_),
    .C(_09241_),
    .D(_09253_),
    .Y(_09254_));
 a31o_1 _13924_ (.A1(_09193_),
    .A2(_09233_),
    .A3(_09241_),
    .B1(_09253_),
    .X(_09255_));
 a2111o_1 _13925_ (.A1(_09254_),
    .A2(_09255_),
    .B1(_09227_),
    .C1(_09244_),
    .D1(_09245_),
    .X(_09256_));
 o311ai_1 _13926_ (.A1(_09227_),
    .A2(_09244_),
    .A3(_09245_),
    .B1(_09254_),
    .C1(_09255_),
    .Y(_09257_));
 a31oi_1 _13927_ (.A1(_09188_),
    .A2(_09256_),
    .A3(_09257_),
    .B1(_09252_),
    .Y(_09258_));
 inv_2 _13928_ (.A(net511),
    .Y(_09259_));
 nand2_1 _13929_ (.A(_09189_),
    .B(_09196_),
    .Y(_09260_));
 o211a_1 _13930_ (.A1(_09189_),
    .A2(_09196_),
    .B1(_09260_),
    .C1(net533),
    .X(_09261_));
 o21ai_1 _13931_ (.A1(_09244_),
    .A2(_09245_),
    .B1(_09227_),
    .Y(_09262_));
 a31oi_4 _13932_ (.A1(_09188_),
    .A2(_09246_),
    .A3(_09262_),
    .B1(_09261_),
    .Y(_09263_));
 inv_2 _13933_ (.A(net508),
    .Y(_09264_));
 or3b_1 _13934_ (.A(_09230_),
    .B(_09242_),
    .C_N(_09237_),
    .X(_09265_));
 and3_1 _13935_ (.A(_09247_),
    .B(_09256_),
    .C(_09265_),
    .X(_09266_));
 nand2_1 _13936_ (.A(_09187_),
    .B(_09232_),
    .Y(_09267_));
 a21o_1 _13937_ (.A1(_09192_),
    .A2(_09231_),
    .B1(_09267_),
    .X(_09268_));
 o31a_1 _13938_ (.A1(net533),
    .A2(_09248_),
    .A3(_09266_),
    .B1(_09268_),
    .X(_09269_));
 o31ai_1 _13939_ (.A1(net533),
    .A2(_09248_),
    .A3(_09266_),
    .B1(_09268_),
    .Y(_09270_));
 nor2_2 _13940_ (.A(net501),
    .B(_09264_),
    .Y(_09271_));
 nor2_1 _13941_ (.A(net501),
    .B(net496),
    .Y(_09272_));
 nand2_2 _13942_ (.A(net500),
    .B(_09271_),
    .Y(_09273_));
 nor2_1 _13943_ (.A(net505),
    .B(_09264_),
    .Y(_09274_));
 a21o_2 _13944_ (.A1(_09234_),
    .A2(_09237_),
    .B1(_09188_),
    .X(_09275_));
 nor2_1 _13945_ (.A(_09234_),
    .B(_09237_),
    .Y(_09276_));
 and2_1 _13946_ (.A(net533),
    .B(_09276_),
    .X(_09277_));
 nand2_4 _13947_ (.A(_09187_),
    .B(_09276_),
    .Y(_09278_));
 nor2_1 _13948_ (.A(_09275_),
    .B(_09276_),
    .Y(_09279_));
 or2_1 _13949_ (.A(_09275_),
    .B(_09276_),
    .X(_09280_));
 and3_1 _13950_ (.A(_09272_),
    .B(_09274_),
    .C(_09275_),
    .X(_09281_));
 and2_1 _13951_ (.A(_09229_),
    .B(_09281_),
    .X(_09282_));
 nor3_1 _13952_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk_before_buf ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.en_ctr ),
    .C(_09282_),
    .Y(_09283_));
 a21oi_1 _13953_ (.A1(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk_before_buf ),
    .A2(\digitop_pav2.sync_inst.inst_clkx.inst_blf.en_ctr ),
    .B1(_09283_),
    .Y(_00576_));
 a21boi_1 _13954_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.pass_t1_i ),
    .A2(_09159_),
    .B1_N(\digitop_pav2.sync_inst.inst_clkx.inst_fm0x.en_fm0x_clk_b ),
    .Y(_00575_));
 nand2_1 _13955_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.dis_blf_fc_b ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.en_blf_fc_b ),
    .Y(_00206_));
 inv_2 _13956_ (.A(_00206_),
    .Y(_00574_));
 a2bb2o_1 _13957_ (.A1_N(net1046),
    .A2_N(_07496_),
    .B1(_07491_),
    .B2(net1038),
    .X(_09284_));
 nor3_1 _13958_ (.A(_07491_),
    .B(_07493_),
    .C(_07547_),
    .Y(_09285_));
 a311o_1 _13959_ (.A1(net1046),
    .A2(_07566_),
    .A3(_09285_),
    .B1(_09284_),
    .C1(_07489_),
    .X(_09286_));
 nor2_1 _13960_ (.A(_07024_),
    .B(_09286_),
    .Y(_09287_));
 or2_1 _13961_ (.A(_07479_),
    .B(_09285_),
    .X(_09288_));
 nand2_1 _13962_ (.A(net1148),
    .B(_07477_),
    .Y(_09289_));
 or4_1 _13963_ (.A(_07491_),
    .B(_07493_),
    .C(_07547_),
    .D(_09289_),
    .X(_09290_));
 nor2_1 _13964_ (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[3] ),
    .B(_09290_),
    .Y(_09291_));
 xor2_1 _13965_ (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[4] ),
    .B(_09291_),
    .X(_09292_));
 a32o_1 _13966_ (.A1(_09287_),
    .A2(_09288_),
    .A3(_09292_),
    .B1(_09286_),
    .B2(\digitop_pav2.access_inst.access_proc0.proc_crc_check[4] ),
    .X(_00370_));
 a31o_1 _13967_ (.A1(net1046),
    .A2(_09288_),
    .A3(_09290_),
    .B1(_09286_),
    .X(_09293_));
 a22o_1 _13968_ (.A1(_09287_),
    .A2(_09291_),
    .B1(_09293_),
    .B2(\digitop_pav2.access_inst.access_proc0.proc_crc_check[3] ),
    .X(_00369_));
 xnor2_1 _13969_ (.A(net1154),
    .B(_07562_),
    .Y(_09294_));
 nand2_1 _13970_ (.A(net1154),
    .B(_07570_),
    .Y(_09295_));
 o21a_1 _13971_ (.A1(_07478_),
    .A2(_07569_),
    .B1(_09295_),
    .X(_09296_));
 nand2_1 _13972_ (.A(net1154),
    .B(_07567_),
    .Y(_09297_));
 a31o_1 _13973_ (.A1(_07548_),
    .A2(_09289_),
    .A3(_09297_),
    .B1(_07493_),
    .X(_09298_));
 a31o_1 _13974_ (.A1(_07479_),
    .A2(_07547_),
    .A3(_09296_),
    .B1(_09298_),
    .X(_09299_));
 nand2_1 _13975_ (.A(\digitop_pav2.access_inst.access_ctrl0.prev_busy ),
    .B(_07578_),
    .Y(_09300_));
 a22o_1 _13976_ (.A1(net1153),
    .A2(_07581_),
    .B1(_09300_),
    .B2(_07477_),
    .X(_09301_));
 nand2_1 _13977_ (.A(_07493_),
    .B(_09301_),
    .Y(_09302_));
 a31o_1 _13978_ (.A1(_07575_),
    .A2(_09299_),
    .A3(_09302_),
    .B1(_09286_),
    .X(_09303_));
 a31o_1 _13979_ (.A1(_07479_),
    .A2(_07491_),
    .A3(_09294_),
    .B1(_09303_),
    .X(_09304_));
 a21bo_1 _13980_ (.A1(net1154),
    .A2(_09286_),
    .B1_N(_09304_),
    .X(_00368_));
 nand2_4 _13981_ (.A(_07511_),
    .B(net912),
    .Y(_09305_));
 a41o_1 _13982_ (.A1(net1234),
    .A2(net818),
    .A3(net965),
    .A4(_09305_),
    .B1(_07616_),
    .X(_09306_));
 a21oi_1 _13983_ (.A1(net965),
    .A2(_07654_),
    .B1(_09306_),
    .Y(_09307_));
 a21bo_1 _13984_ (.A1(net1157),
    .A2(_07631_),
    .B1_N(net202),
    .X(_09308_));
 o21a_1 _13985_ (.A1(net202),
    .A2(_07620_),
    .B1(_09308_),
    .X(_09309_));
 xnor2_1 _13986_ (.A(_07051_),
    .B(_09309_),
    .Y(_09310_));
 a31o_1 _13987_ (.A1(net1157),
    .A2(net1031),
    .A3(_07634_),
    .B1(net1156),
    .X(_09311_));
 o211a_1 _13988_ (.A1(_07513_),
    .A2(_07637_),
    .B1(_07642_),
    .C1(_09311_),
    .X(_09312_));
 a31o_1 _13989_ (.A1(net1157),
    .A2(net1150),
    .A3(net1031),
    .B1(net1156),
    .X(_09313_));
 a31o_1 _13990_ (.A1(_07640_),
    .A2(_07648_),
    .A3(_09313_),
    .B1(_09312_),
    .X(_09314_));
 a22o_1 _13991_ (.A1(net1261),
    .A2(_09310_),
    .B1(_09314_),
    .B2(_07608_),
    .X(_09315_));
 nor2_1 _13992_ (.A(net1156),
    .B(_07620_),
    .Y(_09316_));
 a31o_1 _13993_ (.A1(net1158),
    .A2(net1145),
    .A3(net1032),
    .B1(net1156),
    .X(_09317_));
 a21oi_1 _13994_ (.A1(_07659_),
    .A2(_09317_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.proc_finish0_i ),
    .Y(_09318_));
 o21a_1 _13995_ (.A1(_07738_),
    .A2(_09318_),
    .B1(_07682_),
    .X(_09319_));
 nor2_1 _13996_ (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[5] ),
    .B(_07666_),
    .Y(_09320_));
 or3_1 _13997_ (.A(net1064),
    .B(_07667_),
    .C(_09320_),
    .X(_09321_));
 a31o_1 _13998_ (.A1(net1158),
    .A2(_07568_),
    .A3(net1032),
    .B1(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[5] ),
    .X(_09322_));
 or3b_1 _13999_ (.A(_07672_),
    .B(_07675_),
    .C_N(_09322_),
    .X(_09323_));
 a31o_1 _14000_ (.A1(net1236),
    .A2(_09321_),
    .A3(_09323_),
    .B1(_07511_),
    .X(_09324_));
 a21o_1 _14001_ (.A1(_09319_),
    .A2(_09324_),
    .B1(net1261),
    .X(_09325_));
 or3_1 _14002_ (.A(_07621_),
    .B(_09316_),
    .C(_09319_),
    .X(_09326_));
 o21a_1 _14003_ (.A1(_07621_),
    .A2(_09316_),
    .B1(net1037),
    .X(_09327_));
 a221o_1 _14004_ (.A1(net1071),
    .A2(_07051_),
    .B1(_07627_),
    .B2(_09324_),
    .C1(_09327_),
    .X(_09328_));
 a41o_1 _14005_ (.A1(_07604_),
    .A2(_09325_),
    .A3(_09326_),
    .A4(_09328_),
    .B1(net965),
    .X(_09329_));
 o21ba_1 _14006_ (.A1(_07604_),
    .A2(_09315_),
    .B1_N(_09329_),
    .X(_09330_));
 a21bo_1 _14007_ (.A1(net1073),
    .A2(net965),
    .B1_N(_09307_),
    .X(_09331_));
 o22a_1 _14008_ (.A1(net1156),
    .A2(_09307_),
    .B1(_09330_),
    .B2(_09331_),
    .X(_00367_));
 nor2_1 _14009_ (.A(net1157),
    .B(_07631_),
    .Y(_09332_));
 a21oi_1 _14010_ (.A1(_07559_),
    .A2(net1031),
    .B1(net1158),
    .Y(_09333_));
 or2_1 _14011_ (.A(_07620_),
    .B(_09333_),
    .X(_09334_));
 inv_2 _14012_ (.A(_09334_),
    .Y(_09335_));
 o22a_1 _14013_ (.A1(_09308_),
    .A2(_09332_),
    .B1(_09334_),
    .B2(net201),
    .X(_09336_));
 xor2_1 _14014_ (.A(net1157),
    .B(_07636_),
    .X(_09337_));
 xnor2_1 _14015_ (.A(net1157),
    .B(_07646_),
    .Y(_09338_));
 a22o_1 _14016_ (.A1(_07642_),
    .A2(_09337_),
    .B1(_09338_),
    .B2(_07640_),
    .X(_09339_));
 a2bb2o_1 _14017_ (.A1_N(net1236),
    .A2_N(_09336_),
    .B1(_09339_),
    .B2(_07608_),
    .X(_09340_));
 xor2_1 _14018_ (.A(net1158),
    .B(_07658_),
    .X(_09341_));
 a21oi_1 _14019_ (.A1(_07024_),
    .A2(_09341_),
    .B1(_07738_),
    .Y(_09342_));
 a21oi_1 _14020_ (.A1(net1033),
    .A2(net1032),
    .B1(net1158),
    .Y(_09343_));
 xor2_1 _14021_ (.A(net1158),
    .B(_07671_),
    .X(_09344_));
 o32a_1 _14022_ (.A1(net1064),
    .A2(_07666_),
    .A3(_09343_),
    .B1(_09344_),
    .B2(_07675_),
    .X(_09345_));
 a21oi_1 _14023_ (.A1(net1237),
    .A2(_09345_),
    .B1(_07511_),
    .Y(_09346_));
 o21a_1 _14024_ (.A1(_09342_),
    .A2(_09346_),
    .B1(net1237),
    .X(_09347_));
 nand2_1 _14025_ (.A(_07039_),
    .B(_09334_),
    .Y(_09348_));
 o221a_1 _14026_ (.A1(_07039_),
    .A2(net1158),
    .B1(_07626_),
    .B2(_09346_),
    .C1(_09348_),
    .X(_09349_));
 o211a_1 _14027_ (.A1(_07681_),
    .A2(_09342_),
    .B1(_09335_),
    .C1(_07691_),
    .X(_09350_));
 or4_1 _14028_ (.A(_07603_),
    .B(_09347_),
    .C(_09349_),
    .D(_09350_),
    .X(_09351_));
 o211a_1 _14029_ (.A1(_07604_),
    .A2(_09340_),
    .B1(_09351_),
    .C1(net963),
    .X(_09352_));
 a21bo_1 _14030_ (.A1(net1074),
    .A2(net965),
    .B1_N(_09307_),
    .X(_09353_));
 o22a_1 _14031_ (.A1(net1157),
    .A2(_09307_),
    .B1(_09352_),
    .B2(_09353_),
    .X(_00366_));
 a221o_1 _14032_ (.A1(_07615_),
    .A2(_07653_),
    .B1(_09305_),
    .B2(net964),
    .C1(_07613_),
    .X(_09354_));
 a21o_1 _14033_ (.A1(net964),
    .A2(_07654_),
    .B1(_09354_),
    .X(_09355_));
 nor2_1 _14034_ (.A(net1159),
    .B(_07621_),
    .Y(_09356_));
 or2_1 _14035_ (.A(_07622_),
    .B(_09356_),
    .X(_09357_));
 a21oi_1 _14036_ (.A1(_07512_),
    .A2(_07631_),
    .B1(net1159),
    .Y(_09358_));
 a21o_1 _14037_ (.A1(_07618_),
    .A2(_07631_),
    .B1(_09358_),
    .X(_09359_));
 mux2_1 _14038_ (.A0(_09357_),
    .A1(_09359_),
    .S(net202),
    .X(_09360_));
 inv_2 _14039_ (.A(_09360_),
    .Y(_09361_));
 a31o_1 _14040_ (.A1(_07512_),
    .A2(net1031),
    .A3(_07634_),
    .B1(net1159),
    .X(_09362_));
 and3b_1 _14041_ (.A_N(_07638_),
    .B(_07642_),
    .C(_09362_),
    .X(_09363_));
 or2_1 _14042_ (.A(net1159),
    .B(_07647_),
    .X(_09364_));
 o211a_1 _14043_ (.A1(_07619_),
    .A2(_07646_),
    .B1(_09364_),
    .C1(_07640_),
    .X(_09365_));
 o21a_1 _14044_ (.A1(_09363_),
    .A2(_09365_),
    .B1(_07608_),
    .X(_09366_));
 a211o_1 _14045_ (.A1(net1261),
    .A2(_09361_),
    .B1(_09366_),
    .C1(_07604_),
    .X(_09367_));
 nor2_1 _14046_ (.A(net1159),
    .B(_07672_),
    .Y(_09368_));
 nor2_1 _14047_ (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[6] ),
    .B(_07667_),
    .Y(_09369_));
 a31o_1 _14048_ (.A1(_07577_),
    .A2(net1032),
    .A3(_07618_),
    .B1(_09369_),
    .X(_09370_));
 o32a_1 _14049_ (.A1(_07673_),
    .A2(_07675_),
    .A3(_09368_),
    .B1(_09370_),
    .B2(net1064),
    .X(_09371_));
 or2_1 _14050_ (.A(_07511_),
    .B(_09371_),
    .X(_09372_));
 a22o_1 _14051_ (.A1(\digitop_pav2.access_inst.access_check0.wcnt_check_one ),
    .A2(_07052_),
    .B1(_07628_),
    .B2(_09372_),
    .X(_09373_));
 and2_1 _14052_ (.A(_07052_),
    .B(_07659_),
    .X(_09374_));
 o31a_1 _14053_ (.A1(\digitop_pav2.access_inst.access_ctrl0.proc_finish0_i ),
    .A2(_07660_),
    .A3(_09374_),
    .B1(net1236),
    .X(_09375_));
 a21oi_1 _14054_ (.A1(net1037),
    .A2(_09357_),
    .B1(_09373_),
    .Y(_09376_));
 o22a_1 _14055_ (.A1(net1261),
    .A2(_09372_),
    .B1(_09375_),
    .B2(_07528_),
    .X(_09377_));
 a21oi_1 _14056_ (.A1(net1261),
    .A2(_09357_),
    .B1(_09377_),
    .Y(_09378_));
 o31a_1 _14057_ (.A1(net811),
    .A2(_09376_),
    .A3(_09378_),
    .B1(_07488_),
    .X(_09379_));
 a221o_1 _14058_ (.A1(net1072),
    .A2(net965),
    .B1(_09367_),
    .B2(_09379_),
    .C1(_09355_),
    .X(_09380_));
 a21boi_1 _14059_ (.A1(_07052_),
    .A2(_09355_),
    .B1_N(_09380_),
    .Y(_00365_));
 and2_4 _14060_ (.A(net1481),
    .B(_07055_),
    .X(_09381_));
 mux2_1 _14061_ (.A0(\digitop_pav2.memctrl_inst.addr_to_reram[4] ),
    .A1(net1477),
    .S(_09381_),
    .X(_09382_));
 and2b_2 _14062_ (.A_N(net1481),
    .B(\digitop_pav2.memctrl_inst.busy_ff ),
    .X(_09383_));
 and2_2 _14063_ (.A(net1139),
    .B(net1136),
    .X(_09384_));
 nand2_1 _14064_ (.A(\digitop_pav2.memctrl_inst.addr_to_reram[3] ),
    .B(\digitop_pav2.memctrl_inst.addr_to_reram[4] ),
    .Y(_09385_));
 or4b_1 _14065_ (.A(\digitop_pav2.memctrl_inst.addr_to_reram[1] ),
    .B(_09381_),
    .C(net1027),
    .D_N(\digitop_pav2.memctrl_inst.addr_to_reram[0] ),
    .X(_09386_));
 o22ai_4 _14066_ (.A1(_09381_),
    .A2(_09383_),
    .B1(_09386_),
    .B2(\digitop_pav2.memctrl_inst.addr_to_reram[2] ),
    .Y(_09387_));
 and2b_1 _14067_ (.A_N(_09387_),
    .B(_09382_),
    .X(_09388_));
 nand2b_1 _14068_ (.A_N(_09387_),
    .B(_09382_),
    .Y(_09389_));
 mux2_2 _14069_ (.A0(\digitop_pav2.memctrl_inst.addr_to_reram[1] ),
    .A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[1] ),
    .S(_09381_),
    .X(_09390_));
 mux2_2 _14070_ (.A0(\digitop_pav2.memctrl_inst.addr_to_reram[0] ),
    .A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[0] ),
    .S(_09381_),
    .X(_09391_));
 nor2_1 _14071_ (.A(_09390_),
    .B(_09391_),
    .Y(_09392_));
 inv_2 _14072_ (.A(_09392_),
    .Y(_09393_));
 mux2_2 _14073_ (.A0(\digitop_pav2.memctrl_inst.addr_to_reram[2] ),
    .A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[2] ),
    .S(_09381_),
    .X(_09394_));
 or2_1 _14074_ (.A(_09393_),
    .B(_09394_),
    .X(_09395_));
 or3b_2 _14075_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[0] ),
    .B(net1479),
    .C_N(net1481),
    .X(_09396_));
 o21a_1 _14076_ (.A1(\digitop_pav2.memctrl_inst.addr_to_reram[3] ),
    .A2(_09381_),
    .B1(_09396_),
    .X(_09397_));
 o21ai_4 _14077_ (.A1(\digitop_pav2.memctrl_inst.addr_to_reram[3] ),
    .A2(_09381_),
    .B1(_09396_),
    .Y(_09398_));
 or2_1 _14078_ (.A(_09395_),
    .B(net1025),
    .X(_09399_));
 nor2_1 _14079_ (.A(net957),
    .B(_09399_),
    .Y(net115));
 or3b_1 _14080_ (.A(_09394_),
    .B(_09390_),
    .C_N(_09391_),
    .X(_09400_));
 inv_2 _14081_ (.A(_09400_),
    .Y(_09401_));
 or2_1 _14082_ (.A(net1025),
    .B(_09400_),
    .X(_09402_));
 nor2_1 _14083_ (.A(net957),
    .B(_09402_),
    .Y(net116));
 nand2b_2 _14084_ (.A_N(_09391_),
    .B(_09390_),
    .Y(_09403_));
 or3_1 _14085_ (.A(_09394_),
    .B(net1025),
    .C(_09403_),
    .X(_09404_));
 nor2_1 _14086_ (.A(net957),
    .B(_09404_),
    .Y(net117));
 nand2_1 _14087_ (.A(_09390_),
    .B(_09391_),
    .Y(_09405_));
 nor2_1 _14088_ (.A(_09394_),
    .B(_09405_),
    .Y(_09406_));
 nand2_1 _14089_ (.A(_09398_),
    .B(_09406_),
    .Y(_09407_));
 nor2_1 _14090_ (.A(_09389_),
    .B(_09407_),
    .Y(net118));
 nand2_1 _14091_ (.A(_09392_),
    .B(_09394_),
    .Y(_09408_));
 or2_1 _14092_ (.A(net1025),
    .B(_09408_),
    .X(_09409_));
 nor2_1 _14093_ (.A(net957),
    .B(_09409_),
    .Y(net120));
 nand3b_1 _14094_ (.A_N(_09390_),
    .B(_09391_),
    .C(_09394_),
    .Y(_09410_));
 or2_1 _14095_ (.A(net1025),
    .B(_09410_),
    .X(_09411_));
 nor2_1 _14096_ (.A(net957),
    .B(_09411_),
    .Y(net121));
 and2b_1 _14097_ (.A_N(_09403_),
    .B(_09394_),
    .X(_09412_));
 nand2_1 _14098_ (.A(_09398_),
    .B(_09412_),
    .Y(_09413_));
 nor2_1 _14099_ (.A(net957),
    .B(_09413_),
    .Y(net122));
 and3_1 _14100_ (.A(_09390_),
    .B(_09391_),
    .C(_09394_),
    .X(_09414_));
 and3_1 _14101_ (.A(_09388_),
    .B(_09398_),
    .C(_09414_),
    .X(net123));
 nor2_2 _14102_ (.A(_09382_),
    .B(_09387_),
    .Y(_09415_));
 or2_2 _14103_ (.A(_09382_),
    .B(_09387_),
    .X(_09416_));
 and3_1 _14104_ (.A(_09398_),
    .B(_09414_),
    .C(_09415_),
    .X(net137));
 nor2_1 _14105_ (.A(_09413_),
    .B(net956),
    .Y(net136));
 nor2_1 _14106_ (.A(_09411_),
    .B(net956),
    .Y(net135));
 nor2_1 _14107_ (.A(_09409_),
    .B(net956),
    .Y(net134));
 nor2_1 _14108_ (.A(_09404_),
    .B(net956),
    .Y(net130));
 nor2_1 _14109_ (.A(_09407_),
    .B(_09416_),
    .Y(net133));
 nor2_1 _14110_ (.A(_09399_),
    .B(net956),
    .Y(net108));
 nor2_1 _14111_ (.A(_09402_),
    .B(net956),
    .Y(net119));
 or2_1 _14112_ (.A(_09395_),
    .B(_09398_),
    .X(_09417_));
 nor2_1 _14113_ (.A(net956),
    .B(_09417_),
    .Y(net138));
 and3_1 _14114_ (.A(_09397_),
    .B(_09401_),
    .C(_09415_),
    .X(net139));
 or3_1 _14115_ (.A(_09394_),
    .B(_09398_),
    .C(_09403_),
    .X(_09418_));
 nor2_1 _14116_ (.A(net956),
    .B(_09418_),
    .Y(net109));
 and3_1 _14117_ (.A(_09397_),
    .B(_09406_),
    .C(_09415_),
    .X(net110));
 or2_1 _14118_ (.A(_09398_),
    .B(_09408_),
    .X(_09419_));
 nor2_1 _14119_ (.A(net956),
    .B(_09419_),
    .Y(net111));
 or2_1 _14120_ (.A(_09398_),
    .B(_09410_),
    .X(_09420_));
 nor2_1 _14121_ (.A(net956),
    .B(_09420_),
    .Y(net112));
 and3_1 _14122_ (.A(net1025),
    .B(_09412_),
    .C(_09415_),
    .X(net113));
 and3_1 _14123_ (.A(net1025),
    .B(_09414_),
    .C(_09415_),
    .X(net114));
 nor2_1 _14124_ (.A(_09389_),
    .B(_09417_),
    .Y(net124));
 and4_1 _14125_ (.A(net1477),
    .B(_09381_),
    .C(net1025),
    .D(_09401_),
    .X(net125));
 nor2_1 _14126_ (.A(net957),
    .B(_09418_),
    .Y(net126));
 and3_1 _14127_ (.A(_09388_),
    .B(_09397_),
    .C(_09406_),
    .X(net127));
 nor2_1 _14128_ (.A(net957),
    .B(_09419_),
    .Y(net128));
 nor2_1 _14129_ (.A(net957),
    .B(_09420_),
    .Y(net129));
 and3_1 _14130_ (.A(_09388_),
    .B(net1025),
    .C(_09412_),
    .X(net131));
 and3_1 _14131_ (.A(_09388_),
    .B(net1025),
    .C(_09414_),
    .X(net132));
 nor2_1 _14132_ (.A(_07072_),
    .B(_07931_),
    .Y(_09421_));
 nor2_1 _14133_ (.A(_07958_),
    .B(_09421_),
    .Y(\digitop_pav2.memctrl_inst.n_bit_addr_allow ));
 nor2_1 _14134_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.state[3] ),
    .B(net1488),
    .Y(_09422_));
 or2_1 _14135_ (.A(net1486),
    .B(net1488),
    .X(_09423_));
 nand2_1 _14136_ (.A(net1489),
    .B(net1487),
    .Y(_09424_));
 and3b_1 _14137_ (.A_N(_09424_),
    .B(_07084_),
    .C(net1486),
    .X(_09425_));
 or3_2 _14138_ (.A(net1484),
    .B(_07085_),
    .C(_09424_),
    .X(_09426_));
 nand2_1 _14139_ (.A(net1485),
    .B(\digitop_pav2.testctrl_pav2.inst_mode.state[1] ),
    .Y(_09427_));
 o21a_1 _14140_ (.A1(_09423_),
    .A2(_09427_),
    .B1(_09426_),
    .X(_09428_));
 and2_1 _14141_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.state[3] ),
    .B(net1488),
    .X(_09429_));
 nor2_1 _14142_ (.A(_07085_),
    .B(net1487),
    .Y(_09430_));
 or3_1 _14143_ (.A(_09422_),
    .B(_09427_),
    .C(_09429_),
    .X(_09431_));
 and2_1 _14144_ (.A(net1489),
    .B(net1490),
    .X(_09432_));
 nand2_2 _14145_ (.A(net1489),
    .B(net1490),
    .Y(_09433_));
 a211o_1 _14146_ (.A1(_09422_),
    .A2(_09433_),
    .B1(_09429_),
    .C1(net1485),
    .X(_09434_));
 and4_2 _14147_ (.A(net1489),
    .B(_09428_),
    .C(_09431_),
    .D(_09434_),
    .X(_09435_));
 inv_2 _14148_ (.A(_09435_),
    .Y(_09436_));
 o21a_1 _14149_ (.A1(_09422_),
    .A2(_09435_),
    .B1(net1485),
    .X(_09437_));
 nor2_1 _14150_ (.A(net1485),
    .B(_09423_),
    .Y(_09438_));
 nor2_1 _14151_ (.A(net1489),
    .B(net1490),
    .Y(_09439_));
 and4b_1 _14152_ (.A_N(net1322),
    .B(\digitop_pav2.testctrl_pav2.inst_enter.tm_enter ),
    .C(_09438_),
    .D(_09439_),
    .X(_09440_));
 and3_1 _14153_ (.A(net1502),
    .B(net1504),
    .C(_09440_),
    .X(_09441_));
 nor2_1 _14154_ (.A(_07084_),
    .B(net1486),
    .Y(_09442_));
 nand2_1 _14155_ (.A(net1487),
    .B(_09442_),
    .Y(_09443_));
 nor2_1 _14156_ (.A(net1489),
    .B(_09443_),
    .Y(_09444_));
 nand2_1 _14157_ (.A(net1501),
    .B(net1504),
    .Y(_09445_));
 a311o_1 _14158_ (.A1(net1490),
    .A2(net1501),
    .A3(net1504),
    .B1(_09443_),
    .C1(\digitop_pav2.testctrl_pav2.inst_mode.state[1] ),
    .X(_09446_));
 and2b_1 _14159_ (.A_N(net1504),
    .B(net1502),
    .X(_09447_));
 nand2b_2 _14160_ (.A_N(net1504),
    .B(net1502),
    .Y(_09448_));
 nor2_1 _14161_ (.A(_07084_),
    .B(_07085_),
    .Y(_09449_));
 nand2_1 _14162_ (.A(_09424_),
    .B(_09449_),
    .Y(_09450_));
 nand2_1 _14163_ (.A(_09431_),
    .B(_09450_),
    .Y(_09451_));
 nor2_1 _14164_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.state[1] ),
    .B(net1488),
    .Y(_09452_));
 or2_1 _14165_ (.A(net1489),
    .B(net1487),
    .X(_09453_));
 nor2_1 _14166_ (.A(_09450_),
    .B(_09452_),
    .Y(_09454_));
 a31o_1 _14167_ (.A1(net1490),
    .A2(_09425_),
    .A3(_09447_),
    .B1(_09451_),
    .X(_09455_));
 and2b_1 _14168_ (.A_N(net1489),
    .B(net1491),
    .X(_09456_));
 nand2_1 _14169_ (.A(net1484),
    .B(net1488),
    .Y(_09457_));
 and3_1 _14170_ (.A(net1484),
    .B(net1487),
    .C(_09456_),
    .X(_09458_));
 or4b_2 _14171_ (.A(_09437_),
    .B(_09441_),
    .C(_09455_),
    .D_N(_09446_),
    .X(\digitop_pav2.testctrl_pav2.inst_mode.n_state[4] ));
 inv_2 _14172_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.n_state[4] ),
    .Y(_09459_));
 nor2_1 _14173_ (.A(_09423_),
    .B(_09433_),
    .Y(_09460_));
 and4bb_1 _14174_ (.A_N(net1484),
    .B_N(net1489),
    .C(net1486),
    .D(net1487),
    .X(_09461_));
 a31o_1 _14175_ (.A1(_09432_),
    .A2(_09438_),
    .A3(_09447_),
    .B1(_09461_),
    .X(_09462_));
 and3_2 _14176_ (.A(_07084_),
    .B(_07085_),
    .C(net1487),
    .X(_09463_));
 and3_1 _14177_ (.A(_09432_),
    .B(_09448_),
    .C(_09463_),
    .X(_09464_));
 or3_1 _14178_ (.A(net1484),
    .B(_07085_),
    .C(net1487),
    .X(_09465_));
 or2_1 _14179_ (.A(_09433_),
    .B(_09465_),
    .X(_09466_));
 inv_2 _14180_ (.A(_09466_),
    .Y(_09467_));
 a31o_1 _14181_ (.A1(net1501),
    .A2(net1504),
    .A3(_09467_),
    .B1(_09464_),
    .X(_09468_));
 and3_1 _14182_ (.A(net1487),
    .B(_09439_),
    .C(_09449_),
    .X(_09469_));
 or4_1 _14183_ (.A(_07084_),
    .B(net1487),
    .C(_09433_),
    .D(_09448_),
    .X(_09470_));
 a221o_1 _14184_ (.A1(net1486),
    .A2(_09458_),
    .B1(_09463_),
    .B2(_09433_),
    .C1(_09469_),
    .X(_09471_));
 or3b_1 _14185_ (.A(_09444_),
    .B(_09462_),
    .C_N(_09470_),
    .X(_09472_));
 a211o_1 _14186_ (.A1(net1501),
    .A2(_09440_),
    .B1(_09468_),
    .C1(_09472_),
    .X(_09473_));
 a21oi_1 _14187_ (.A1(net1490),
    .A2(_09447_),
    .B1(_09426_),
    .Y(_09474_));
 and2b_1 _14188_ (.A_N(net1490),
    .B(net1489),
    .X(_09475_));
 nand2b_1 _14189_ (.A_N(_09443_),
    .B(_09475_),
    .Y(_09476_));
 nor2_1 _14190_ (.A(_09433_),
    .B(_09443_),
    .Y(_09477_));
 nand2_1 _14191_ (.A(_09448_),
    .B(_09477_),
    .Y(_09478_));
 or4bb_1 _14192_ (.A(_09435_),
    .B(_09474_),
    .C_N(_09476_),
    .D_N(_09478_),
    .X(_09479_));
 o32a_2 _14193_ (.A1(_09471_),
    .A2(_09473_),
    .A3(_09479_),
    .B1(_09436_),
    .B2(net1484),
    .X(\digitop_pav2.testctrl_pav2.inst_mode.n_state[2] ));
 a22o_1 _14194_ (.A1(_09449_),
    .A2(_09452_),
    .B1(_09477_),
    .B2(_09447_),
    .X(_09480_));
 and3_1 _14195_ (.A(net1484),
    .B(_09430_),
    .C(_09432_),
    .X(_09481_));
 nor2_1 _14196_ (.A(_09432_),
    .B(_09465_),
    .Y(_09482_));
 or4_1 _14197_ (.A(_09441_),
    .B(_09474_),
    .C(_09481_),
    .D(_09482_),
    .X(_09483_));
 a32o_1 _14198_ (.A1(net1501),
    .A2(_09432_),
    .A3(_09463_),
    .B1(_09458_),
    .B2(net1486),
    .X(_09484_));
 a41o_1 _14199_ (.A1(_07085_),
    .A2(net1501),
    .A3(net1504),
    .A4(_09458_),
    .B1(_09462_),
    .X(_09485_));
 and3_1 _14200_ (.A(net1484),
    .B(_09430_),
    .C(_09475_),
    .X(_09486_));
 nor2_1 _14201_ (.A(_09469_),
    .B(_09486_),
    .Y(_09487_));
 o21ai_1 _14202_ (.A1(net1501),
    .A2(_09466_),
    .B1(_09487_),
    .Y(_09488_));
 a211o_1 _14203_ (.A1(_09445_),
    .A2(_09484_),
    .B1(_09485_),
    .C1(_09488_),
    .X(_09489_));
 or3_1 _14204_ (.A(_09480_),
    .B(_09483_),
    .C(_09489_),
    .X(_09490_));
 nor2_1 _14205_ (.A(_09474_),
    .B(_09485_),
    .Y(_09491_));
 a21oi_2 _14206_ (.A1(net1486),
    .A2(_09435_),
    .B1(_09490_),
    .Y(_09492_));
 inv_2 _14207_ (.A(_09492_),
    .Y(\digitop_pav2.testctrl_pav2.inst_mode.n_state[3] ));
 a22o_1 _14208_ (.A1(_09445_),
    .A2(_09467_),
    .B1(_09481_),
    .B2(_09448_),
    .X(_09493_));
 or3_1 _14209_ (.A(net1490),
    .B(_09423_),
    .C(_09427_),
    .X(_09494_));
 o211a_1 _14210_ (.A1(net1484),
    .A2(_09423_),
    .B1(_09456_),
    .C1(_09457_),
    .X(_09495_));
 a31o_1 _14211_ (.A1(net1504),
    .A2(_09438_),
    .A3(_09456_),
    .B1(_09447_),
    .X(_09496_));
 o22a_1 _14212_ (.A1(_09448_),
    .A2(_09495_),
    .B1(_09496_),
    .B2(_09460_),
    .X(_09497_));
 a21bo_1 _14213_ (.A1(net1501),
    .A2(_09458_),
    .B1_N(_09494_),
    .X(_09498_));
 o21a_1 _14214_ (.A1(_09430_),
    .A2(_09463_),
    .B1(_09475_),
    .X(_09499_));
 or4_1 _14215_ (.A(_09464_),
    .B(_09493_),
    .C(_09498_),
    .D(_09499_),
    .X(_09500_));
 nor4_1 _14216_ (.A(_09441_),
    .B(_09479_),
    .C(_09497_),
    .D(_09500_),
    .Y(_09501_));
 inv_2 _14217_ (.A(net1309),
    .Y(\digitop_pav2.testctrl_pav2.inst_mode.n_state[1] ));
 a21oi_1 _14218_ (.A1(net67),
    .A2(_09440_),
    .B1(_09458_),
    .Y(_09502_));
 nor2_1 _14219_ (.A(net1502),
    .B(_09502_),
    .Y(_09503_));
 and2b_1 _14220_ (.A_N(net1501),
    .B(net1504),
    .X(_09504_));
 o31a_1 _14221_ (.A1(_09460_),
    .A2(_09495_),
    .A3(_09503_),
    .B1(_09448_),
    .X(_09505_));
 and3b_1 _14222_ (.A_N(_09504_),
    .B(_09456_),
    .C(_09438_),
    .X(_09506_));
 a311o_1 _14223_ (.A1(net1490),
    .A2(_09425_),
    .A3(_09448_),
    .B1(_09464_),
    .C1(_09506_),
    .X(_09507_));
 or4b_1 _14224_ (.A(_07084_),
    .B(net1491),
    .C(net1486),
    .D_N(_09424_),
    .X(_09508_));
 a211o_1 _14225_ (.A1(net1485),
    .A2(_09453_),
    .B1(_09422_),
    .C1(net1491),
    .X(_09509_));
 a31o_1 _14226_ (.A1(_09487_),
    .A2(_09508_),
    .A3(_09509_),
    .B1(_09448_),
    .X(_09510_));
 o21ai_1 _14227_ (.A1(_09448_),
    .A2(_09476_),
    .B1(_09478_),
    .Y(_09511_));
 or4b_1 _14228_ (.A(_09493_),
    .B(_09511_),
    .C(_09507_),
    .D_N(_09510_),
    .X(_09512_));
 a211o_1 _14229_ (.A1(net1490),
    .A2(_09435_),
    .B1(_09505_),
    .C1(_09512_),
    .X(\digitop_pav2.testctrl_pav2.inst_mode.n_state[0] ));
 a31o_1 _14230_ (.A1(\digitop_pav2.access_inst.access_ctrl0.dt_acc_done_o ),
    .A2(\digitop_pav2.access_inst.access_ctrl0.state[15] ),
    .A3(net1191),
    .B1(\digitop_pav2.access_inst.access_ctrl0.state[1] ),
    .X(_00025_));
 a22o_1 _14231_ (.A1(net1248),
    .A2(\digitop_pav2.ack_inst.state_ff[0] ),
    .B1(_08872_),
    .B2(\digitop_pav2.ack_inst.state_ff[2] ),
    .X(_00041_));
 or3b_1 _14232_ (.A(\digitop_pav2.ack_inst.rcnt_ff[1] ),
    .B(net1234),
    .C_N(_08510_),
    .X(_09513_));
 a22o_1 _14233_ (.A1(\digitop_pav2.ack_inst.nvm_ack_rd_stb_o ),
    .A2(net1248),
    .B1(_09513_),
    .B2(\digitop_pav2.ack_inst.state_ff[1] ),
    .X(_00040_));
 nand2_1 _14234_ (.A(\digitop_pav2.access_inst.access_ctrl0.tx_dt_finish_i ),
    .B(net1191),
    .Y(_09514_));
 nor2_1 _14235_ (.A(net1208),
    .B(net818),
    .Y(_09515_));
 inv_2 _14236_ (.A(_09515_),
    .Y(_09516_));
 or2_1 _14237_ (.A(\digitop_pav2.access_inst.access_ctrl0.replay_nok ),
    .B(net1260),
    .X(_09517_));
 a32o_1 _14238_ (.A1(_08472_),
    .A2(_09515_),
    .A3(_09517_),
    .B1(_09514_),
    .B2(net1142),
    .X(_00031_));
 mux2_1 _14239_ (.A0(_07555_),
    .A1(\digitop_pav2.access_inst.access_ctrl0.state[24] ),
    .S(_07960_),
    .X(_00030_));
 nor2_1 _14240_ (.A(net1235),
    .B(_07104_),
    .Y(_09518_));
 and3_1 _14241_ (.A(\digitop_pav2.access_inst.access_check0.pc_lock_check_sync_o ),
    .B(net1238),
    .C(net1699),
    .X(_09519_));
 nand2b_1 _14242_ (.A_N(\digitop_pav2.access_inst.access_check0.fg_i[4] ),
    .B(\digitop_pav2.access_inst.access_check0.permalock_tid_i ),
    .Y(_09520_));
 a31oi_2 _14243_ (.A1(net1260),
    .A2(net811),
    .A3(_09520_),
    .B1(\digitop_pav2.access_inst.access_check0.lock_error_o ),
    .Y(_09521_));
 a31o_1 _14244_ (.A1(net1260),
    .A2(net811),
    .A3(_09520_),
    .B1(\digitop_pav2.access_inst.access_check0.lock_error_o ),
    .X(_09522_));
 nor2_1 _14245_ (.A(\digitop_pav2.access_inst.access_check0.pc_invalid_o ),
    .B(_09522_),
    .Y(_09523_));
 nor2_1 _14246_ (.A(_07033_),
    .B(_07576_),
    .Y(_09524_));
 and3_1 _14247_ (.A(net1152),
    .B(net1191),
    .C(_07395_),
    .X(_09525_));
 nor2_1 _14248_ (.A(_07034_),
    .B(_07987_),
    .Y(_09526_));
 a32o_1 _14249_ (.A1(net1046),
    .A2(net1145),
    .A3(net1190),
    .B1(_07960_),
    .B2(\digitop_pav2.access_inst.access_ctrl0.state[23] ),
    .X(_09527_));
 a31o_1 _14250_ (.A1(net1067),
    .A2(\digitop_pav2.access_inst.access_ctrl0.state[11] ),
    .A3(_07959_),
    .B1(_09527_),
    .X(_09528_));
 a41o_1 _14251_ (.A1(net1650),
    .A2(net1700),
    .A3(_07970_),
    .A4(_09526_),
    .B1(_09528_),
    .X(_09529_));
 a31o_1 _14252_ (.A1(net1318),
    .A2(_09524_),
    .A3(_09525_),
    .B1(_09529_),
    .X(_09530_));
 a31o_1 _14253_ (.A1(_09518_),
    .A2(_09519_),
    .A3(_09523_),
    .B1(_09530_),
    .X(_00029_));
 a32o_1 _14254_ (.A1(net1258),
    .A2(net1143),
    .A3(_07334_),
    .B1(net1205),
    .B2(\digitop_pav2.access_inst.access_ctrl0.state[22] ),
    .X(_00028_));
 a22o_1 _14255_ (.A1(\digitop_pav2.access_inst.access_ctrl0.ld_dt_stb ),
    .A2(net1205),
    .B1(_07959_),
    .B2(\digitop_pav2.access_inst.access_ctrl0.state[14] ),
    .X(_00027_));
 nand2_1 _14256_ (.A(net1194),
    .B(net819),
    .Y(_09531_));
 a32o_1 _14257_ (.A1(\digitop_pav2.access_inst.access_ctrl0.rx_par0_i ),
    .A2(\digitop_pav2.access_inst.access_ctrl0.state[13] ),
    .A3(_07396_),
    .B1(_09531_),
    .B2(\digitop_pav2.access_inst.access_ctrl0.state[20] ),
    .X(_00026_));
 o211a_1 _14258_ (.A1(net1067),
    .A2(net1318),
    .B1(_07575_),
    .C1(_07033_),
    .X(_09532_));
 o2111a_1 _14259_ (.A1(_07396_),
    .A2(_09532_),
    .B1(_08470_),
    .C1(net1152),
    .D1(net1191),
    .X(_09533_));
 a2bb2o_1 _14260_ (.A1_N(\digitop_pav2.access_inst.access_ctrl0.nvm_busy_i ),
    .A2_N(_07554_),
    .B1(_09516_),
    .B2(net1143),
    .X(_09534_));
 a211o_1 _14261_ (.A1(\digitop_pav2.access_inst.access_ctrl0.state[5] ),
    .A2(net1191),
    .B1(_09533_),
    .C1(_09534_),
    .X(_00024_));
 mux2_1 _14262_ (.A0(\digitop_pav2.access_inst.access_ctrl0.state[24] ),
    .A1(\digitop_pav2.access_inst.access_ctrl0.state[18] ),
    .S(_07960_),
    .X(_00023_));
 a22o_1 _14263_ (.A1(\digitop_pav2.access_inst.access_check0.wr_lock_ck_i ),
    .A2(net1206),
    .B1(_07959_),
    .B2(\digitop_pav2.access_inst.access_ctrl0.state[2] ),
    .X(_00021_));
 o21a_1 _14264_ (.A1(_07022_),
    .A2(_09531_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.state[17] ),
    .X(_09535_));
 nand2_1 _14265_ (.A(\digitop_pav2.access_inst.access_ctrl0.rx_par0_i ),
    .B(net1194),
    .Y(_09536_));
 a41o_1 _14266_ (.A1(\digitop_pav2.access_inst.access_ctrl0.rx_par0_i ),
    .A2(\digitop_pav2.access_inst.access_ctrl0.state[13] ),
    .A3(net1194),
    .A4(_07395_),
    .B1(_09535_),
    .X(_00022_));
 a22o_4 _14267_ (.A1(net1180),
    .A2(net578),
    .B1(net536),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_m[1] ),
    .X(_09537_));
 a22o_2 _14268_ (.A1(net1179),
    .A2(net578),
    .B1(net536),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_m[0] ),
    .X(_09538_));
 inv_2 _14269_ (.A(_09538_),
    .Y(_09539_));
 nor2_1 _14270_ (.A(_09537_),
    .B(_09538_),
    .Y(_09540_));
 or2_1 _14271_ (.A(_09537_),
    .B(_09538_),
    .X(_09541_));
 and2_1 _14272_ (.A(_08520_),
    .B(net531),
    .X(_09542_));
 or3b_1 _14273_ (.A(_09539_),
    .B(_09537_),
    .C_N(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[0] ),
    .X(_09543_));
 inv_2 _14274_ (.A(_09543_),
    .Y(_09544_));
 and3_1 _14275_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[2] ),
    .B(_09537_),
    .C(_09539_),
    .X(_09545_));
 nand2_1 _14276_ (.A(_09537_),
    .B(_09538_),
    .Y(_09546_));
 and3_1 _14277_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[6] ),
    .B(_09537_),
    .C(_09538_),
    .X(_09547_));
 nor4_1 _14278_ (.A(_09542_),
    .B(_09544_),
    .C(_09545_),
    .D(_09547_),
    .Y(_09548_));
 or3_1 _14279_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_trext ),
    .B(_07256_),
    .C(_07270_),
    .X(_09549_));
 o31a_1 _14280_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[5] ),
    .A2(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[12] ),
    .A3(_07327_),
    .B1(_09549_),
    .X(_09550_));
 a221o_4 _14281_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[3] ),
    .A2(net578),
    .B1(net536),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_trext ),
    .C1(_09550_),
    .X(_09551_));
 inv_2 _14282_ (.A(_09551_),
    .Y(_09552_));
 nand2_1 _14283_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[1] ),
    .B(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[0] ),
    .Y(_09553_));
 or3_1 _14284_ (.A(_07122_),
    .B(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[3] ),
    .C(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[2] ),
    .X(_09554_));
 o21ai_1 _14285_ (.A1(_09553_),
    .A2(_09554_),
    .B1(_09551_),
    .Y(_09555_));
 nor2_1 _14286_ (.A(net188),
    .B(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[3] ),
    .Y(_09556_));
 nand2_1 _14287_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[2] ),
    .B(_09556_),
    .Y(_09557_));
 nor2_1 _14288_ (.A(_09553_),
    .B(_09557_),
    .Y(_09558_));
 o21a_1 _14289_ (.A1(_09551_),
    .A2(_09558_),
    .B1(_09555_),
    .X(_09559_));
 or3_1 _14290_ (.A(net188),
    .B(_07124_),
    .C(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[2] ),
    .X(_09560_));
 or2_1 _14291_ (.A(_09553_),
    .B(_09560_),
    .X(_09561_));
 nor2_1 _14292_ (.A(_09551_),
    .B(_09561_),
    .Y(_09562_));
 and3_1 _14293_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[1] ),
    .B(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[0] ),
    .C(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[2] ),
    .X(_09563_));
 a41o_1 _14294_ (.A1(net188),
    .A2(_07124_),
    .A3(_09551_),
    .A4(_09563_),
    .B1(net531),
    .X(_09564_));
 o22a_1 _14295_ (.A1(net530),
    .A2(_09559_),
    .B1(_09562_),
    .B2(_09564_),
    .X(_09565_));
 nand2_1 _14296_ (.A(_09548_),
    .B(_09565_),
    .Y(\digitop_pav2.fm0miller_inst.fm0x_ctrl.n_data_valid ));
 nor2_1 _14297_ (.A(net1399),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.piex_dt_rx_done ),
    .Y(_00169_));
 or2_2 _14298_ (.A(\digitop_pav2.memctrl_inst.ctr[0] ),
    .B(\digitop_pav2.memctrl_inst.ctr[1] ),
    .X(_09566_));
 or3_1 _14299_ (.A(\digitop_pav2.memctrl_inst.ctr[2] ),
    .B(\digitop_pav2.memctrl_inst.ctr[3] ),
    .C(\digitop_pav2.memctrl_inst.ctr[4] ),
    .X(_09567_));
 or2_1 _14300_ (.A(\digitop_pav2.memctrl_inst.ctr[5] ),
    .B(_09567_),
    .X(_09568_));
 or2_1 _14301_ (.A(_09566_),
    .B(_09568_),
    .X(_09569_));
 or2_1 _14302_ (.A(\digitop_pav2.memctrl_inst.ctr[6] ),
    .B(_09569_),
    .X(_09570_));
 nor2_1 _14303_ (.A(\digitop_pav2.memctrl_inst.ctr[7] ),
    .B(_09570_),
    .Y(_09571_));
 o31a_1 _14304_ (.A1(\digitop_pav2.memctrl_inst.ctr[7] ),
    .A2(_07139_),
    .A3(_09570_),
    .B1(\digitop_pav2.memctrl_inst.state[3] ),
    .X(\digitop_pav2.memctrl_inst.n_read ));
 nor2_1 _14305_ (.A(\digitop_pav2.func_rr_prog ),
    .B(\digitop_pav2.func_rr_erase ),
    .Y(_09572_));
 and3b_1 _14306_ (.A_N(_09572_),
    .B(_09571_),
    .C(\digitop_pav2.memctrl_inst.state[4] ),
    .X(\digitop_pav2.memctrl_inst.n_state[2] ));
 or2_1 _14307_ (.A(\digitop_pav2.pie_inst.fsm.dif_pos_fix[0] ),
    .B(\digitop_pav2.pie_inst.fsm.past_ctr[1] ),
    .X(_09573_));
 or2_1 _14308_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[2] ),
    .B(_09573_),
    .X(_09574_));
 nand2_1 _14309_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[2] ),
    .B(_09573_),
    .Y(_09575_));
 nand2_2 _14310_ (.A(_09574_),
    .B(_09575_),
    .Y(_09576_));
 inv_2 _14311_ (.A(_09576_),
    .Y(\digitop_pav2.pie_inst.fsm.dif_pos_fix[2] ));
 or2_4 _14312_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[3] ),
    .B(_09574_),
    .X(_09577_));
 inv_2 _14313_ (.A(_09577_),
    .Y(_09578_));
 or3_1 _14314_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[4] ),
    .B(\digitop_pav2.pie_inst.fsm.past_ctr[5] ),
    .C(_09577_),
    .X(_09579_));
 or2_1 _14315_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[6] ),
    .B(_09579_),
    .X(_09580_));
 xnor2_1 _14316_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[7] ),
    .B(_09580_),
    .Y(_09581_));
 inv_2 _14317_ (.A(net494),
    .Y(\digitop_pav2.pie_inst.fsm.dif_pos_fix[7] ));
 nand2_1 _14318_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[3] ),
    .B(_09574_),
    .Y(_09582_));
 nand2_2 _14319_ (.A(_09577_),
    .B(_09582_),
    .Y(_09583_));
 inv_2 _14320_ (.A(_09583_),
    .Y(\digitop_pav2.pie_inst.fsm.dif_pos_fix[3] ));
 or3_2 _14321_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[7] ),
    .B(\digitop_pav2.pie_inst.fsm.past_ctr[8] ),
    .C(_09580_),
    .X(_09584_));
 xnor2_4 _14322_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[9] ),
    .B(_09584_),
    .Y(_09585_));
 inv_2 _14323_ (.A(_09585_),
    .Y(\digitop_pav2.pie_inst.fsm.dif_pos_fix[9] ));
 nand2_1 _14324_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[6] ),
    .B(_09579_),
    .Y(_09586_));
 nand2_1 _14325_ (.A(_09580_),
    .B(_09586_),
    .Y(_09587_));
 inv_2 _14326_ (.A(net493),
    .Y(\digitop_pav2.pie_inst.fsm.dif_pos_fix[6] ));
 o21ai_1 _14327_ (.A1(\digitop_pav2.pie_inst.fsm.past_ctr[4] ),
    .A2(_09577_),
    .B1(\digitop_pav2.pie_inst.fsm.past_ctr[5] ),
    .Y(_09588_));
 nand2_1 _14328_ (.A(_09579_),
    .B(_09588_),
    .Y(_09589_));
 inv_2 _14329_ (.A(net495),
    .Y(\digitop_pav2.pie_inst.fsm.dif_pos_fix[5] ));
 or2_1 _14330_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[1] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[2] ),
    .X(_09590_));
 nor4_1 _14331_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[0] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[3] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[4] ),
    .D(_09590_),
    .Y(_09591_));
 or4_4 _14332_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[0] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[3] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[4] ),
    .D(_09590_),
    .X(_09592_));
 and4_1 _14333_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[4] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[5] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[7] ),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[6] ),
    .X(_09593_));
 and3_1 _14334_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[0] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[1] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[2] ),
    .X(_09594_));
 and3_1 _14335_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[3] ),
    .B(_09593_),
    .C(_09594_),
    .X(_09595_));
 and4_1 _14336_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[9] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[8] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[11] ),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[10] ),
    .X(_09596_));
 and4_1 _14337_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[13] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[12] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[15] ),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[14] ),
    .X(_09597_));
 and3_2 _14338_ (.A(_09595_),
    .B(_09596_),
    .C(_09597_),
    .X(_09598_));
 nand3_2 _14339_ (.A(_09595_),
    .B(_09596_),
    .C(_09597_),
    .Y(_09599_));
 a21o_1 _14340_ (.A1(_09592_),
    .A2(_09598_),
    .B1(_07152_),
    .X(_09600_));
 nor2_1 _14341_ (.A(_07151_),
    .B(_09592_),
    .Y(_09601_));
 nand2_1 _14342_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_end_i ),
    .B(net1466),
    .Y(_09602_));
 a22o_1 _14343_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[2] ),
    .A2(_09600_),
    .B1(_09601_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[7] ),
    .X(_00117_));
 and4_1 _14344_ (.A(net1480),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[2] ),
    .C(net1466),
    .D(_09598_),
    .X(_09603_));
 a21o_1 _14345_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[6] ),
    .A2(_09602_),
    .B1(_09603_),
    .X(_00121_));
 or4_1 _14346_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[4] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[5] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[7] ),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[6] ),
    .X(_09604_));
 or4_1 _14347_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[0] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[1] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[2] ),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[3] ),
    .X(_09605_));
 or4_1 _14348_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[9] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[8] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[11] ),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[10] ),
    .X(_09606_));
 or4_1 _14349_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[13] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[12] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[15] ),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[14] ),
    .X(_09607_));
 or3_1 _14350_ (.A(_09604_),
    .B(_09605_),
    .C(_09607_),
    .X(_09608_));
 nor2_4 _14351_ (.A(_09606_),
    .B(_09608_),
    .Y(_09609_));
 a21o_1 _14352_ (.A1(_09592_),
    .A2(_09609_),
    .B1(_07152_),
    .X(_09610_));
 a22o_1 _14353_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[5] ),
    .A2(_09601_),
    .B1(_09610_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[3] ),
    .X(_00118_));
 a22o_1 _14354_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[6] ),
    .A2(_09601_),
    .B1(_09610_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[4] ),
    .X(_00119_));
 and4_1 _14355_ (.A(net1480),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[3] ),
    .C(net1466),
    .D(_09609_),
    .X(_09611_));
 a21o_1 _14356_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[7] ),
    .A2(_09602_),
    .B1(_09611_),
    .X(_00122_));
 nand2_1 _14357_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[2] ),
    .B(_09599_),
    .Y(_09612_));
 nor2_1 _14358_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[3] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[4] ),
    .Y(_09613_));
 o21ai_1 _14359_ (.A1(_09609_),
    .A2(_09613_),
    .B1(_09612_),
    .Y(_09614_));
 a21o_1 _14360_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rd_end_i ),
    .A2(_09614_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[1] ),
    .X(_00116_));
 a22o_1 _14361_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.form_end ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[0] ),
    .B1(_09602_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[5] ),
    .X(_00120_));
 a41o_1 _14362_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rd_end_i ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[4] ),
    .A3(net1466),
    .A4(_09609_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[8] ),
    .X(_00123_));
 nand2_1 _14363_ (.A(net1481),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[0] ),
    .Y(_09615_));
 mux2_1 _14364_ (.A0(net1501),
    .A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[2] ),
    .S(_09615_),
    .X(_00124_));
 mux2_1 _14365_ (.A0(_09504_),
    .A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[3] ),
    .S(_09615_),
    .X(_00125_));
 a22o_1 _14366_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_end_i ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[5] ),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[3] ),
    .B2(_07152_),
    .X(_00106_));
 a22o_1 _14367_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_end_i ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[7] ),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[2] ),
    .B2(_07152_),
    .X(_00105_));
 nand2_1 _14368_ (.A(net1480),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[2] ),
    .Y(_09616_));
 or4_1 _14369_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[2] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[5] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[6] ),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[7] ),
    .X(_09617_));
 or4_1 _14370_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[0] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[1] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[3] ),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[4] ),
    .X(_09618_));
 nor4_1 _14371_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[9] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[8] ),
    .C(_09617_),
    .D(_09618_),
    .Y(_09619_));
 or4_1 _14372_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[9] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[8] ),
    .C(_09617_),
    .D(_09618_),
    .X(_09620_));
 or3b_1 _14373_ (.A(_09599_),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[3] ),
    .C_N(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.read_after_prog_ok ),
    .X(_09621_));
 nor2_1 _14374_ (.A(_09616_),
    .B(_09621_),
    .Y(_09622_));
 a211o_1 _14375_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[8] ),
    .A2(net1465),
    .B1(_09622_),
    .C1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_form_end ),
    .X(_09623_));
 or4_1 _14376_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[0] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[4] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[5] ),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[6] ),
    .X(_09624_));
 or4_1 _14377_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[1] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[2] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[3] ),
    .D(_09624_),
    .X(_09625_));
 or4_4 _14378_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[7] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[9] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[8] ),
    .D(_09625_),
    .X(_09626_));
 inv_2 _14379_ (.A(_09626_),
    .Y(_09627_));
 a31o_1 _14380_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[1] ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[0] ),
    .A3(_09627_),
    .B1(_09623_),
    .X(_00104_));
 or2_2 _14381_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.int_wr_stb ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_stb ),
    .X(_09628_));
 nor3_1 _14382_ (.A(_07055_),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.int_rd_stb ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rd_stb ),
    .Y(_09629_));
 nor3_1 _14383_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.int_rd_stb ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rd_stb ),
    .C(_09628_),
    .Y(_09630_));
 or3_2 _14384_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.int_rd_stb ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rd_stb ),
    .C(_09628_),
    .X(_09631_));
 or3_2 _14385_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[0] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[1] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[2] ),
    .X(_09632_));
 or3_2 _14386_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[3] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[4] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[5] ),
    .X(_09633_));
 nor2_4 _14387_ (.A(_09632_),
    .B(_09633_),
    .Y(_09634_));
 or2_2 _14388_ (.A(_09632_),
    .B(_09633_),
    .X(_09635_));
 or4_2 _14389_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[0] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[1] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[3] ),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[2] ),
    .X(_09636_));
 inv_2 _14390_ (.A(_09636_),
    .Y(_09637_));
 a21o_1 _14391_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[1] ),
    .A2(_09637_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[4] ),
    .X(_09638_));
 a22o_1 _14392_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[0] ),
    .A2(_09630_),
    .B1(_09634_),
    .B2(_09638_),
    .X(_00112_));
 mux2_1 _14393_ (.A0(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[1] ),
    .A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[2] ),
    .S(_09634_),
    .X(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_state[2] ));
 a22o_1 _14394_ (.A1(_09628_),
    .A2(_09629_),
    .B1(_09635_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[2] ),
    .X(_09639_));
 a31o_1 _14395_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[1] ),
    .A2(_09634_),
    .A3(_09636_),
    .B1(_09639_),
    .X(_00113_));
 a21oi_2 _14396_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.rr_read ),
    .A2(_09634_),
    .B1(_07156_),
    .Y(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_read ));
 o21a_1 _14397_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.int_rd_stb ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rd_stb ),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[0] ),
    .X(_09640_));
 or2_1 _14398_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_read ),
    .B(_09640_),
    .X(_00114_));
 and3_1 _14399_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.rr_read ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[3] ),
    .C(_09634_),
    .X(_09641_));
 a21o_1 _14400_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[4] ),
    .A2(_09635_),
    .B1(_09641_),
    .X(_00115_));
 or3_1 _14401_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[1] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[2] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[3] ),
    .X(_09642_));
 nor3_1 _14402_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[0] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[4] ),
    .C(_09642_),
    .Y(_09643_));
 nand2_1 _14403_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_end_i ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[4] ),
    .Y(_09644_));
 a32o_1 _14404_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_end_i ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[4] ),
    .A3(_09643_),
    .B1(_09620_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[8] ),
    .X(_00111_));
 and2_1 _14405_ (.A(net1480),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[3] ),
    .X(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_int_wr_bit ));
 a21o_1 _14406_ (.A1(_07151_),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[7] ),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_int_wr_bit ),
    .X(_00110_));
 a32o_1 _14407_ (.A1(net1480),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[2] ),
    .A3(_09621_),
    .B1(_09620_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[6] ),
    .X(_00109_));
 and3b_1 _14408_ (.A_N(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[1] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[0] ),
    .C(_09627_),
    .X(_09645_));
 a21o_1 _14409_ (.A1(_07151_),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[5] ),
    .B1(_09645_),
    .X(_00108_));
 and2_1 _14410_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[6] ),
    .B(net1465),
    .X(_09646_));
 nand2_1 _14411_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_end_i ),
    .B(_09643_),
    .Y(_09647_));
 a21o_1 _14412_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[4] ),
    .A2(_09647_),
    .B1(_09646_),
    .X(_00107_));
 o21ai_1 _14413_ (.A1(\digitop_pav2.pie_inst.fsm.past_ctr[7] ),
    .A2(_09580_),
    .B1(\digitop_pav2.pie_inst.fsm.past_ctr[8] ),
    .Y(_09648_));
 nand2_1 _14414_ (.A(_09584_),
    .B(_09648_),
    .Y(_09649_));
 inv_2 _14415_ (.A(net491),
    .Y(\digitop_pav2.pie_inst.fsm.dif_pos_fix[8] ));
 or3_1 _14416_ (.A(\digitop_pav2.sec_inst.shift_out.st[2] ),
    .B(\digitop_pav2.sec_inst.shift_out.st[4] ),
    .C(_08503_),
    .X(_09650_));
 a31o_1 _14417_ (.A1(\digitop_pav2.sec_inst.shift_out.st[5] ),
    .A2(_08505_),
    .A3(_08507_),
    .B1(\digitop_pav2.sec_inst.shift_out.st[7] ),
    .X(_00103_));
 o21a_1 _14418_ (.A1(net707),
    .A2(_08505_),
    .B1(_09650_),
    .X(_00102_));
 a211o_1 _14419_ (.A1(_07064_),
    .A2(net701),
    .B1(_08504_),
    .C1(net709),
    .X(_09651_));
 o21a_1 _14420_ (.A1(\digitop_pav2.sec_inst.shift_out.st[5] ),
    .A2(_08505_),
    .B1(_09651_),
    .X(_00101_));
 mux2_1 _14421_ (.A0(_08506_),
    .A1(net709),
    .S(_08504_),
    .X(_00100_));
 nor2_1 _14422_ (.A(\digitop_pav2.sec_inst.ld_mem.st[1] ),
    .B(_09165_),
    .Y(_09652_));
 a21boi_1 _14423_ (.A1(\digitop_pav2.sec_inst.ld_mem.st[3] ),
    .A2(net1635),
    .B1_N(_09652_),
    .Y(_09653_));
 o21ba_1 _14424_ (.A1(\digitop_pav2.sec_inst.ld_mem.st[1] ),
    .A2(\digitop_pav2.sec_inst.ld_mem.st[0] ),
    .B1_N(net1636),
    .X(_09654_));
 or2_1 _14425_ (.A(net715),
    .B(_07108_),
    .X(_09655_));
 or2_1 _14426_ (.A(\digitop_pav2.sec_inst.ld_mem.wctr[0] ),
    .B(\digitop_pav2.sec_inst.ld_mem.wctr[1] ),
    .X(_09656_));
 a21oi_1 _14427_ (.A1(\digitop_pav2.sec_inst.ld_mem.wctr[3] ),
    .A2(_09655_),
    .B1(_09656_),
    .Y(_09657_));
 xnor2_1 _14428_ (.A(\digitop_pav2.sec_inst.ld_mem.wctr[2] ),
    .B(_07852_),
    .Y(_09658_));
 o211ai_1 _14429_ (.A1(\digitop_pav2.sec_inst.ld_mem.wctr[3] ),
    .A2(_09655_),
    .B1(_09657_),
    .C1(_09658_),
    .Y(_09659_));
 or2_1 _14430_ (.A(\digitop_pav2.sec_inst.ld_mem.st[1] ),
    .B(net1636),
    .X(_09660_));
 nand2_1 _14431_ (.A(\digitop_pav2.sec_inst.ld_mem.st[2] ),
    .B(_09660_),
    .Y(_09661_));
 a31o_1 _14432_ (.A1(\digitop_pav2.sec_inst.ld_mem.st[2] ),
    .A2(_09659_),
    .A3(_09660_),
    .B1(_09654_),
    .X(_00098_));
 nor2_1 _14433_ (.A(_09659_),
    .B(_09661_),
    .Y(_00099_));
 a21o_1 _14434_ (.A1(\digitop_pav2.access_inst.access_ctrl0.tx_dt_finish_i ),
    .A2(net1142),
    .B1(\digitop_pav2.access_inst.access_ctrl0.state[22] ),
    .X(_09662_));
 a22o_1 _14435_ (.A1(\digitop_pav2.access_inst.access_ctrl0.state[15] ),
    .A2(_08466_),
    .B1(_09662_),
    .B2(net1191),
    .X(_09663_));
 a41o_1 _14436_ (.A1(_07037_),
    .A2(net1238),
    .A3(_08472_),
    .A4(_09515_),
    .B1(_09663_),
    .X(_00020_));
 and2_1 _14437_ (.A(net970),
    .B(\digitop_pav2.proc_ctrl_inst.ebv.state[0] ),
    .X(_09664_));
 a22o_1 _14438_ (.A1(_07111_),
    .A2(\digitop_pav2.proc_ctrl_inst.ebv.state[8] ),
    .B1(_09664_),
    .B2(net1299),
    .X(_00097_));
 nor2_1 _14439_ (.A(net499),
    .B(net516),
    .Y(_09665_));
 nor2_1 _14440_ (.A(net503),
    .B(net511),
    .Y(_09666_));
 nor2_1 _14441_ (.A(net509),
    .B(net499),
    .Y(_09667_));
 xnor2_2 _14442_ (.A(_09264_),
    .B(net499),
    .Y(_09668_));
 nor2_1 _14443_ (.A(net523),
    .B(net510),
    .Y(_09669_));
 a21oi_2 _14444_ (.A1(_09223_),
    .A2(_09224_),
    .B1(_09220_),
    .Y(_09670_));
 or3_2 _14445_ (.A(_09185_),
    .B(_09188_),
    .C(_09204_),
    .X(_09671_));
 o31ai_4 _14446_ (.A1(net533),
    .A2(_09225_),
    .A3(_09670_),
    .B1(_09671_),
    .Y(_09672_));
 o31a_1 _14447_ (.A1(net533),
    .A2(_09225_),
    .A3(_09670_),
    .B1(_09671_),
    .X(_09673_));
 nor2_2 _14448_ (.A(net508),
    .B(net513),
    .Y(_09674_));
 xnor2_2 _14449_ (.A(_09229_),
    .B(net510),
    .Y(_09675_));
 a21o_1 _14450_ (.A1(_09674_),
    .A2(_09675_),
    .B1(_09669_),
    .X(_09676_));
 a21o_1 _14451_ (.A1(_09668_),
    .A2(_09676_),
    .B1(_09667_),
    .X(_09677_));
 nor2_1 _14452_ (.A(net506),
    .B(net502),
    .Y(_09678_));
 nor2_1 _14453_ (.A(_09666_),
    .B(_09678_),
    .Y(_09679_));
 a21o_2 _14454_ (.A1(_09677_),
    .A2(_09679_),
    .B1(_09666_),
    .X(_09680_));
 nand2_1 _14455_ (.A(net499),
    .B(net516),
    .Y(_09681_));
 and2b_1 _14456_ (.A_N(_09665_),
    .B(_09681_),
    .X(_09682_));
 a21oi_2 _14457_ (.A1(_09680_),
    .A2(_09681_),
    .B1(_09665_),
    .Y(_09683_));
 nor2_2 _14458_ (.A(net506),
    .B(net520),
    .Y(_09684_));
 inv_2 _14459_ (.A(_09684_),
    .Y(_09685_));
 xnor2_4 _14460_ (.A(_09683_),
    .B(_09684_),
    .Y(_09686_));
 and2_1 _14461_ (.A(\digitop_pav2.pie_inst.fsm.pivot[7] ),
    .B(_09686_),
    .X(_09687_));
 xnor2_4 _14462_ (.A(_09680_),
    .B(_09682_),
    .Y(_09688_));
 or2_1 _14463_ (.A(net1300),
    .B(_09688_),
    .X(_09689_));
 xnor2_1 _14464_ (.A(net1300),
    .B(_09688_),
    .Y(_09690_));
 xnor2_2 _14465_ (.A(_09677_),
    .B(_09679_),
    .Y(_09691_));
 nand2_1 _14466_ (.A(\digitop_pav2.pie_inst.fsm.pivot[5] ),
    .B(_09691_),
    .Y(_09692_));
 or2_1 _14467_ (.A(\digitop_pav2.pie_inst.fsm.pivot[5] ),
    .B(_09691_),
    .X(_09693_));
 xnor2_2 _14468_ (.A(_09668_),
    .B(_09676_),
    .Y(_09694_));
 inv_2 _14469_ (.A(_09694_),
    .Y(_09695_));
 and2_1 _14470_ (.A(\digitop_pav2.pie_inst.fsm.pivot[4] ),
    .B(_09694_),
    .X(_09696_));
 or2_1 _14471_ (.A(\digitop_pav2.pie_inst.fsm.pivot[4] ),
    .B(_09694_),
    .X(_09697_));
 and2b_1 _14472_ (.A_N(_09696_),
    .B(_09697_),
    .X(_09698_));
 xor2_2 _14473_ (.A(_09674_),
    .B(_09675_),
    .X(_09699_));
 xnor2_1 _14474_ (.A(_09674_),
    .B(_09675_),
    .Y(_09700_));
 and2_1 _14475_ (.A(net1301),
    .B(_09700_),
    .X(_09701_));
 nand2_1 _14476_ (.A(net1301),
    .B(_09700_),
    .Y(_09702_));
 nor2_1 _14477_ (.A(net1301),
    .B(_09700_),
    .Y(_09703_));
 xnor2_4 _14478_ (.A(_09263_),
    .B(_09672_),
    .Y(_09704_));
 xnor2_2 _14479_ (.A(net508),
    .B(net512),
    .Y(_09705_));
 and2_1 _14480_ (.A(\digitop_pav2.pie_inst.fsm.pivot[2] ),
    .B(_09705_),
    .X(_09706_));
 xnor2_2 _14481_ (.A(\digitop_pav2.pie_inst.fsm.pivot[2] ),
    .B(_09704_),
    .Y(_09707_));
 and2_1 _14482_ (.A(\digitop_pav2.pie_inst.fsm.pivot[1] ),
    .B(net523),
    .X(_09708_));
 or2_1 _14483_ (.A(\digitop_pav2.pie_inst.fsm.pivot[1] ),
    .B(net523),
    .X(_09709_));
 xnor2_1 _14484_ (.A(\digitop_pav2.pie_inst.fsm.pivot[1] ),
    .B(net523),
    .Y(_09710_));
 nor2_1 _14485_ (.A(\digitop_pav2.pie_inst.fsm.pivot[0] ),
    .B(net512),
    .Y(_09711_));
 nor2_1 _14486_ (.A(_09710_),
    .B(_09711_),
    .Y(_09712_));
 or2_1 _14487_ (.A(_09708_),
    .B(_09712_),
    .X(_09713_));
 a21oi_1 _14488_ (.A1(_09707_),
    .A2(_09713_),
    .B1(_09706_),
    .Y(_09714_));
 a21oi_1 _14489_ (.A1(_09702_),
    .A2(_09714_),
    .B1(_09703_),
    .Y(_09715_));
 a21o_1 _14490_ (.A1(_09697_),
    .A2(_09715_),
    .B1(_09696_),
    .X(_09716_));
 nand2_1 _14491_ (.A(_09693_),
    .B(_09716_),
    .Y(_09717_));
 a21oi_1 _14492_ (.A1(_09692_),
    .A2(_09717_),
    .B1(_09690_),
    .Y(_09718_));
 a21oi_1 _14493_ (.A1(net1300),
    .A2(_09688_),
    .B1(_09718_),
    .Y(_09719_));
 o211ai_1 _14494_ (.A1(net498),
    .A2(_09680_),
    .B1(_09685_),
    .C1(net518),
    .Y(_09720_));
 a31o_1 _14495_ (.A1(net497),
    .A2(_09680_),
    .A3(_09685_),
    .B1(net518),
    .X(_09721_));
 nand2_1 _14496_ (.A(_09720_),
    .B(_09721_),
    .Y(_09722_));
 nand2_2 _14497_ (.A(\digitop_pav2.pie_inst.fsm.pivot[8] ),
    .B(_09722_),
    .Y(_09723_));
 nor2_1 _14498_ (.A(\digitop_pav2.pie_inst.fsm.pivot[7] ),
    .B(_09686_),
    .Y(_09724_));
 o21ba_1 _14499_ (.A1(_09719_),
    .A2(_09724_),
    .B1_N(_09687_),
    .X(_09725_));
 or2_2 _14500_ (.A(_09723_),
    .B(_09725_),
    .X(_09726_));
 inv_2 _14501_ (.A(_09726_),
    .Y(_09727_));
 xnor2_1 _14502_ (.A(net510),
    .B(net518),
    .Y(_09728_));
 nor2_1 _14503_ (.A(_09250_),
    .B(net509),
    .Y(_09729_));
 nor2_1 _14504_ (.A(net522),
    .B(net499),
    .Y(_09730_));
 nor2_1 _14505_ (.A(_09229_),
    .B(net497),
    .Y(_09731_));
 nor2_1 _14506_ (.A(_09730_),
    .B(_09731_),
    .Y(_09732_));
 nor2_1 _14507_ (.A(net510),
    .B(net512),
    .Y(_09733_));
 and2_1 _14508_ (.A(_09732_),
    .B(_09733_),
    .X(_09734_));
 nor2_1 _14509_ (.A(_09274_),
    .B(_09729_),
    .Y(_09735_));
 o21a_1 _14510_ (.A1(_09730_),
    .A2(_09734_),
    .B1(_09735_),
    .X(_09736_));
 o21ai_1 _14511_ (.A1(_09729_),
    .A2(_09736_),
    .B1(_09728_),
    .Y(_09737_));
 o21ai_1 _14512_ (.A1(net510),
    .A2(net516),
    .B1(_09737_),
    .Y(_09738_));
 o21ai_1 _14513_ (.A1(net497),
    .A2(net521),
    .B1(_09738_),
    .Y(_09739_));
 nor2_1 _14514_ (.A(net503),
    .B(_09739_),
    .Y(_09740_));
 xnor2_1 _14515_ (.A(net516),
    .B(_09740_),
    .Y(_09741_));
 nand2_1 _14516_ (.A(net478),
    .B(_09741_),
    .Y(_09742_));
 nor2_1 _14517_ (.A(\digitop_pav2.pie_inst.fsm.pivot[8] ),
    .B(_09722_),
    .Y(_09743_));
 nor2_1 _14518_ (.A(_07149_),
    .B(_09672_),
    .Y(_09744_));
 o221a_1 _14519_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[2] ),
    .A2(_09705_),
    .B1(_09708_),
    .B2(_09744_),
    .C1(_09709_),
    .X(_09745_));
 a211oi_1 _14520_ (.A1(net1301),
    .A2(_09700_),
    .B1(_09706_),
    .C1(_09745_),
    .Y(_09746_));
 a2bb2o_1 _14521_ (.A1_N(_09703_),
    .A2_N(_09746_),
    .B1(\digitop_pav2.pie_inst.fsm.pivot[4] ),
    .B2(_09694_),
    .X(_09747_));
 a22o_1 _14522_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[5] ),
    .A2(_09691_),
    .B1(_09697_),
    .B2(_09747_),
    .X(_09748_));
 a22o_1 _14523_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[6] ),
    .A2(_09688_),
    .B1(_09693_),
    .B2(_09748_),
    .X(_09749_));
 a22oi_1 _14524_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[7] ),
    .A2(_09686_),
    .B1(_09689_),
    .B2(_09749_),
    .Y(_09750_));
 nor2_1 _14525_ (.A(_09687_),
    .B(_09724_),
    .Y(_09751_));
 o31ai_1 _14526_ (.A1(_09724_),
    .A2(_09743_),
    .A3(_09750_),
    .B1(_09723_),
    .Y(_09752_));
 o31a_2 _14527_ (.A1(_09724_),
    .A2(_09743_),
    .A3(_09750_),
    .B1(_09723_),
    .X(_09753_));
 nand2_1 _14528_ (.A(_09719_),
    .B(_09751_),
    .Y(_09754_));
 or2_1 _14529_ (.A(_09719_),
    .B(_09751_),
    .X(_09755_));
 a21o_1 _14530_ (.A1(_09754_),
    .A2(_09755_),
    .B1(_09753_),
    .X(_09756_));
 inv_2 _14531_ (.A(net476),
    .Y(_09757_));
 and2_1 _14532_ (.A(net503),
    .B(_09739_),
    .X(_09758_));
 nor2_1 _14533_ (.A(_09740_),
    .B(_09758_),
    .Y(_09759_));
 o22ai_1 _14534_ (.A1(_09726_),
    .A2(_09741_),
    .B1(net476),
    .B2(_09759_),
    .Y(_09760_));
 and3_1 _14535_ (.A(_09690_),
    .B(_09692_),
    .C(_09717_),
    .X(_09761_));
 or3_1 _14536_ (.A(_09718_),
    .B(_09753_),
    .C(_09761_),
    .X(_09762_));
 inv_2 _14537_ (.A(net486),
    .Y(_09763_));
 or3_1 _14538_ (.A(net497),
    .B(net521),
    .C(_09738_),
    .X(_09764_));
 and2_1 _14539_ (.A(_09739_),
    .B(_09764_),
    .X(_09765_));
 nor2_1 _14540_ (.A(net486),
    .B(_09765_),
    .Y(_09766_));
 nand2_1 _14541_ (.A(_09692_),
    .B(_09693_),
    .Y(_09767_));
 xnor2_2 _14542_ (.A(_09716_),
    .B(_09767_),
    .Y(_09768_));
 nand2_2 _14543_ (.A(net490),
    .B(_09768_),
    .Y(_09769_));
 inv_2 _14544_ (.A(net484),
    .Y(_09770_));
 or3_1 _14545_ (.A(_09728_),
    .B(_09729_),
    .C(_09736_),
    .X(_09771_));
 and2_1 _14546_ (.A(_09737_),
    .B(_09771_),
    .X(_09772_));
 nor2_1 _14547_ (.A(_09769_),
    .B(_09772_),
    .Y(_09773_));
 nand2_1 _14548_ (.A(net484),
    .B(_09772_),
    .Y(_09774_));
 and2b_1 _14549_ (.A_N(_09773_),
    .B(_09774_),
    .X(_09775_));
 xor2_1 _14550_ (.A(_09698_),
    .B(_09715_),
    .X(_09776_));
 nand2_1 _14551_ (.A(net489),
    .B(_09776_),
    .Y(_09777_));
 nor3_1 _14552_ (.A(_09730_),
    .B(_09734_),
    .C(_09735_),
    .Y(_09778_));
 nor2_1 _14553_ (.A(_09736_),
    .B(_09778_),
    .Y(_09779_));
 nor2_1 _14554_ (.A(net483),
    .B(_09779_),
    .Y(_09780_));
 and2_1 _14555_ (.A(net483),
    .B(_09779_),
    .X(_09781_));
 nor2_1 _14556_ (.A(_09780_),
    .B(_09781_),
    .Y(_09782_));
 nor2_1 _14557_ (.A(_09701_),
    .B(_09703_),
    .Y(_09783_));
 xnor2_1 _14558_ (.A(_09714_),
    .B(_09783_),
    .Y(_09784_));
 and2_2 _14559_ (.A(net489),
    .B(_09784_),
    .X(_09785_));
 nand2_1 _14560_ (.A(net489),
    .B(_09784_),
    .Y(_09786_));
 nor2_1 _14561_ (.A(_09732_),
    .B(_09733_),
    .Y(_09787_));
 or2_1 _14562_ (.A(_09734_),
    .B(_09787_),
    .X(_09788_));
 xnor2_1 _14563_ (.A(_09785_),
    .B(_09788_),
    .Y(_09789_));
 inv_2 _14564_ (.A(_09789_),
    .Y(_09790_));
 xor2_2 _14565_ (.A(_09707_),
    .B(_09713_),
    .X(_09791_));
 nand2_1 _14566_ (.A(net487),
    .B(_09791_),
    .Y(_09792_));
 nor2_1 _14567_ (.A(net502),
    .B(net514),
    .Y(_09793_));
 nor2_1 _14568_ (.A(_09733_),
    .B(_09793_),
    .Y(_09794_));
 nor2_1 _14569_ (.A(net479),
    .B(_09794_),
    .Y(_09795_));
 nand2_1 _14570_ (.A(net479),
    .B(_09794_),
    .Y(_09796_));
 and2_1 _14571_ (.A(_09710_),
    .B(_09711_),
    .X(_09797_));
 nor2_1 _14572_ (.A(_09712_),
    .B(_09797_),
    .Y(_09798_));
 and2_1 _14573_ (.A(net487),
    .B(net492),
    .X(_09799_));
 and3_1 _14574_ (.A(net509),
    .B(net488),
    .C(_09798_),
    .X(_09800_));
 or2_1 _14575_ (.A(_09711_),
    .B(_09744_),
    .X(_09801_));
 and2_1 _14576_ (.A(net487),
    .B(_09801_),
    .X(_09802_));
 or3b_2 _14577_ (.A(_09229_),
    .B(_09753_),
    .C_N(_09801_),
    .X(_09803_));
 a21o_2 _14578_ (.A1(net489),
    .A2(_09801_),
    .B1(net523),
    .X(_09804_));
 and3_1 _14579_ (.A(net513),
    .B(_09803_),
    .C(_09804_),
    .X(_09805_));
 a21bo_2 _14580_ (.A1(net512),
    .A2(_09804_),
    .B1_N(_09803_),
    .X(_09806_));
 a21o_1 _14581_ (.A1(net488),
    .A2(_09798_),
    .B1(net509),
    .X(_09807_));
 and2b_1 _14582_ (.A_N(_09800_),
    .B(_09807_),
    .X(_09808_));
 a21o_1 _14583_ (.A1(_09806_),
    .A2(_09807_),
    .B1(_09800_),
    .X(_09809_));
 a211o_1 _14584_ (.A1(_09806_),
    .A2(_09807_),
    .B1(_09795_),
    .C1(_09800_),
    .X(_09810_));
 nand2_1 _14585_ (.A(_09796_),
    .B(_09810_),
    .Y(_09811_));
 a32o_1 _14586_ (.A1(_09790_),
    .A2(_09796_),
    .A3(_09810_),
    .B1(_09788_),
    .B2(_09785_),
    .X(_09812_));
 a21o_1 _14587_ (.A1(_09782_),
    .A2(_09812_),
    .B1(_09780_),
    .X(_09813_));
 a21o_1 _14588_ (.A1(_09774_),
    .A2(_09813_),
    .B1(_09773_),
    .X(_09814_));
 nand2_1 _14589_ (.A(net486),
    .B(_09765_),
    .Y(_09815_));
 nand2b_1 _14590_ (.A_N(_09766_),
    .B(_09815_),
    .Y(_09816_));
 a21o_1 _14591_ (.A1(_09814_),
    .A2(_09815_),
    .B1(_09766_),
    .X(_09817_));
 nand2_1 _14592_ (.A(net477),
    .B(_09759_),
    .Y(_09818_));
 inv_2 _14593_ (.A(_09818_),
    .Y(_09819_));
 a21o_1 _14594_ (.A1(_09817_),
    .A2(_09818_),
    .B1(_09760_),
    .X(_09820_));
 xnor2_2 _14595_ (.A(net518),
    .B(net478),
    .Y(_09821_));
 xnor2_1 _14596_ (.A(net503),
    .B(net477),
    .Y(_09822_));
 o21ai_1 _14597_ (.A1(net498),
    .A2(net486),
    .B1(_09822_),
    .Y(_09823_));
 nor2_1 _14598_ (.A(net499),
    .B(_09763_),
    .Y(_09824_));
 nor2_1 _14599_ (.A(_09264_),
    .B(net483),
    .Y(_09825_));
 xnor2_1 _14600_ (.A(net509),
    .B(net483),
    .Y(_09826_));
 and3_1 _14601_ (.A(net523),
    .B(net489),
    .C(_09784_),
    .X(_09827_));
 a21o_1 _14602_ (.A1(net489),
    .A2(_09791_),
    .B1(net512),
    .X(_09828_));
 a21o_1 _14603_ (.A1(net489),
    .A2(_09784_),
    .B1(net523),
    .X(_09829_));
 nand2b_1 _14604_ (.A_N(_09827_),
    .B(_09829_),
    .Y(_09830_));
 a21o_1 _14605_ (.A1(_09828_),
    .A2(_09829_),
    .B1(_09827_),
    .X(_09831_));
 a21oi_1 _14606_ (.A1(_09826_),
    .A2(_09831_),
    .B1(_09825_),
    .Y(_09832_));
 a221o_1 _14607_ (.A1(net510),
    .A2(_09770_),
    .B1(_09826_),
    .B2(_09831_),
    .C1(_09825_),
    .X(_09833_));
 o21ai_1 _14608_ (.A1(net510),
    .A2(_09770_),
    .B1(_09833_),
    .Y(_09834_));
 or3_1 _14609_ (.A(_09823_),
    .B(_09824_),
    .C(_09834_),
    .X(_09835_));
 a211o_1 _14610_ (.A1(net506),
    .A2(net477),
    .B1(net486),
    .C1(net498),
    .X(_09836_));
 o211a_1 _14611_ (.A1(net506),
    .A2(net477),
    .B1(_09835_),
    .C1(_09836_),
    .X(_09837_));
 xnor2_1 _14612_ (.A(net510),
    .B(_09769_),
    .Y(_09838_));
 o32ai_4 _14613_ (.A1(net518),
    .A2(_09723_),
    .A3(_09725_),
    .B1(_09821_),
    .B2(_09837_),
    .Y(_09839_));
 o211ai_1 _14614_ (.A1(_09822_),
    .A2(_09824_),
    .B1(_09834_),
    .C1(_09823_),
    .Y(_09840_));
 xnor2_1 _14615_ (.A(_09832_),
    .B(_09838_),
    .Y(_09841_));
 xor2_1 _14616_ (.A(_09826_),
    .B(_09831_),
    .X(_09842_));
 nor2_1 _14617_ (.A(net511),
    .B(net508),
    .Y(_09843_));
 a21oi_1 _14618_ (.A1(_09263_),
    .A2(_09802_),
    .B1(net510),
    .Y(_09844_));
 a21oi_1 _14619_ (.A1(_09271_),
    .A2(_09802_),
    .B1(_09799_),
    .Y(_09845_));
 or2_1 _14620_ (.A(_09844_),
    .B(_09845_),
    .X(_09846_));
 or2_1 _14621_ (.A(net497),
    .B(_09846_),
    .X(_09847_));
 o22a_1 _14622_ (.A1(net514),
    .A2(net479),
    .B1(_09846_),
    .B2(net497),
    .X(_09848_));
 and2_1 _14623_ (.A(net497),
    .B(_09846_),
    .X(_09849_));
 xnor2_1 _14624_ (.A(_09828_),
    .B(_09830_),
    .Y(_09850_));
 nor2_1 _14625_ (.A(_09250_),
    .B(_09850_),
    .Y(_09851_));
 a211oi_1 _14626_ (.A1(_09828_),
    .A2(_09848_),
    .B1(_09849_),
    .C1(_09851_),
    .Y(_09852_));
 a221o_1 _14627_ (.A1(net516),
    .A2(_09842_),
    .B1(_09850_),
    .B2(_09250_),
    .C1(_09852_),
    .X(_09853_));
 nor2_1 _14628_ (.A(_09278_),
    .B(_09770_),
    .Y(_09854_));
 nand2_2 _14629_ (.A(net520),
    .B(net484),
    .Y(_09855_));
 or2_1 _14630_ (.A(net516),
    .B(_09842_),
    .X(_09856_));
 a32o_1 _14631_ (.A1(_09853_),
    .A2(_09855_),
    .A3(_09856_),
    .B1(_09841_),
    .B2(_09278_),
    .X(_09857_));
 xor2_1 _14632_ (.A(_09821_),
    .B(_09837_),
    .X(_09858_));
 a211o_1 _14633_ (.A1(_09835_),
    .A2(_09840_),
    .B1(_09857_),
    .C1(_09858_),
    .X(_09859_));
 a22o_1 _14634_ (.A1(_09742_),
    .A2(_09820_),
    .B1(_09839_),
    .B2(_09859_),
    .X(_09860_));
 nor2_1 _14635_ (.A(net504),
    .B(net519),
    .Y(_09861_));
 nand2_1 _14636_ (.A(net504),
    .B(net519),
    .Y(_09862_));
 nor2_1 _14637_ (.A(_09250_),
    .B(net500),
    .Y(_09863_));
 nor2_1 _14638_ (.A(net511),
    .B(net500),
    .Y(_09864_));
 or2_1 _14639_ (.A(_09271_),
    .B(_09843_),
    .X(_09865_));
 a21o_1 _14640_ (.A1(net508),
    .A2(net513),
    .B1(net522),
    .X(_09866_));
 nor2_1 _14641_ (.A(_09865_),
    .B(_09866_),
    .Y(_09867_));
 nor2_1 _14642_ (.A(_09272_),
    .B(_09864_),
    .Y(_09868_));
 o21ai_1 _14643_ (.A1(_09843_),
    .A2(_09867_),
    .B1(_09868_),
    .Y(_09869_));
 nand2b_2 _14644_ (.A_N(_09864_),
    .B(_09869_),
    .Y(_09870_));
 nor2_1 _14645_ (.A(net504),
    .B(net498),
    .Y(_09871_));
 nor2_2 _14646_ (.A(_09863_),
    .B(_09871_),
    .Y(_09872_));
 a21oi_4 _14647_ (.A1(_09870_),
    .A2(_09872_),
    .B1(_09863_),
    .Y(_09873_));
 o21a_1 _14648_ (.A1(_09861_),
    .A2(_09873_),
    .B1(_09862_),
    .X(_09874_));
 nor2_1 _14649_ (.A(_09275_),
    .B(_09874_),
    .Y(_09875_));
 or2_1 _14650_ (.A(net520),
    .B(_09875_),
    .X(_09876_));
 nor2_2 _14651_ (.A(net478),
    .B(_09876_),
    .Y(_09877_));
 nor2_1 _14652_ (.A(_09275_),
    .B(_09875_),
    .Y(_09878_));
 and2b_1 _14653_ (.A_N(_09874_),
    .B(_09275_),
    .X(_09879_));
 or2_1 _14654_ (.A(_09878_),
    .B(_09879_),
    .X(_09880_));
 nor2_1 _14655_ (.A(net504),
    .B(_09878_),
    .Y(_09881_));
 nor2_1 _14656_ (.A(_09879_),
    .B(_09881_),
    .Y(_09882_));
 and2b_1 _14657_ (.A_N(_09861_),
    .B(_09862_),
    .X(_09883_));
 xor2_4 _14658_ (.A(_09873_),
    .B(_09883_),
    .X(_09884_));
 xor2_2 _14659_ (.A(_09870_),
    .B(_09872_),
    .X(_09885_));
 nand2_1 _14660_ (.A(net501),
    .B(_09885_),
    .Y(_09886_));
 xnor2_1 _14661_ (.A(net511),
    .B(_09885_),
    .Y(_09887_));
 or3_1 _14662_ (.A(_09843_),
    .B(_09867_),
    .C(_09868_),
    .X(_09888_));
 and2_1 _14663_ (.A(_09869_),
    .B(_09888_),
    .X(_09889_));
 and2_1 _14664_ (.A(_09264_),
    .B(_09889_),
    .X(_09890_));
 nor2_1 _14665_ (.A(_09264_),
    .B(_09889_),
    .Y(_09891_));
 or2_1 _14666_ (.A(_09890_),
    .B(_09891_),
    .X(_09892_));
 and2_1 _14667_ (.A(_09865_),
    .B(_09866_),
    .X(_09893_));
 nor2_1 _14668_ (.A(_09867_),
    .B(_09893_),
    .Y(_09894_));
 a22oi_1 _14669_ (.A1(net511),
    .A2(_09674_),
    .B1(_09894_),
    .B2(_09229_),
    .Y(_09895_));
 nor2_1 _14670_ (.A(_09892_),
    .B(_09895_),
    .Y(_09896_));
 o21ai_1 _14671_ (.A1(_09890_),
    .A2(_09896_),
    .B1(_09887_),
    .Y(_09897_));
 xnor2_1 _14672_ (.A(net500),
    .B(_09884_),
    .Y(_09898_));
 a21o_1 _14673_ (.A1(_09886_),
    .A2(_09897_),
    .B1(_09898_),
    .X(_09899_));
 o21a_1 _14674_ (.A1(net500),
    .A2(_09884_),
    .B1(_09899_),
    .X(_09900_));
 o21ba_1 _14675_ (.A1(_09881_),
    .A2(_09900_),
    .B1_N(_09879_),
    .X(_09901_));
 and2b_1 _14676_ (.A_N(_09901_),
    .B(_09878_),
    .X(_09902_));
 and2b_1 _14677_ (.A_N(_09878_),
    .B(_09901_),
    .X(_09903_));
 nor2_1 _14678_ (.A(_09902_),
    .B(_09903_),
    .Y(_09904_));
 nor2_1 _14679_ (.A(net476),
    .B(_09904_),
    .Y(_09905_));
 xnor2_1 _14680_ (.A(_09882_),
    .B(_09900_),
    .Y(_09906_));
 and2_1 _14681_ (.A(net485),
    .B(_09906_),
    .X(_09907_));
 nor2_1 _14682_ (.A(net485),
    .B(_09906_),
    .Y(_09908_));
 nand3_1 _14683_ (.A(_09886_),
    .B(_09897_),
    .C(_09898_),
    .Y(_09909_));
 and2_1 _14684_ (.A(_09899_),
    .B(_09909_),
    .X(_09910_));
 xnor2_1 _14685_ (.A(_09770_),
    .B(_09910_),
    .Y(_09911_));
 or3_1 _14686_ (.A(_09887_),
    .B(_09890_),
    .C(_09896_),
    .X(_09912_));
 and2_1 _14687_ (.A(_09897_),
    .B(_09912_),
    .X(_09913_));
 nor2_1 _14688_ (.A(net482),
    .B(_09913_),
    .Y(_09914_));
 nand2_1 _14689_ (.A(net482),
    .B(_09913_),
    .Y(_09915_));
 and2_1 _14690_ (.A(_09892_),
    .B(_09895_),
    .X(_09916_));
 nor2_1 _14691_ (.A(_09896_),
    .B(_09916_),
    .Y(_09917_));
 nor2_1 _14692_ (.A(net481),
    .B(_09917_),
    .Y(_09918_));
 nand2_1 _14693_ (.A(net481),
    .B(_09917_),
    .Y(_09919_));
 nand2b_1 _14694_ (.A_N(_09918_),
    .B(_09919_),
    .Y(_09920_));
 nand2_1 _14695_ (.A(net522),
    .B(net508),
    .Y(_09921_));
 nand2_1 _14696_ (.A(net513),
    .B(_09921_),
    .Y(_09922_));
 xnor2_1 _14697_ (.A(net501),
    .B(_09922_),
    .Y(_09923_));
 or2_1 _14698_ (.A(net479),
    .B(_09923_),
    .X(_09924_));
 nand2_1 _14699_ (.A(net479),
    .B(_09923_),
    .Y(_09925_));
 nor2_1 _14700_ (.A(_09229_),
    .B(net514),
    .Y(_09926_));
 o21ai_2 _14701_ (.A1(net522),
    .A2(_09705_),
    .B1(_09921_),
    .Y(_09927_));
 a21o_1 _14702_ (.A1(net513),
    .A2(_09927_),
    .B1(_09674_),
    .X(_09928_));
 and3_1 _14703_ (.A(net488),
    .B(net492),
    .C(_09928_),
    .X(_09929_));
 nand2_1 _14704_ (.A(net522),
    .B(net514),
    .Y(_09930_));
 nand2_1 _14705_ (.A(_09804_),
    .B(_09930_),
    .Y(_09931_));
 a21o_1 _14706_ (.A1(net488),
    .A2(_09798_),
    .B1(_09928_),
    .X(_09932_));
 nand2b_1 _14707_ (.A_N(_09929_),
    .B(_09932_),
    .Y(_09933_));
 or2_1 _14708_ (.A(_09931_),
    .B(_09933_),
    .X(_09934_));
 a31oi_2 _14709_ (.A1(_09804_),
    .A2(_09930_),
    .A3(_09932_),
    .B1(_09929_),
    .Y(_09935_));
 nand2_1 _14710_ (.A(_09924_),
    .B(_09935_),
    .Y(_09936_));
 nand2_1 _14711_ (.A(_09925_),
    .B(_09936_),
    .Y(_09937_));
 a31o_1 _14712_ (.A1(_09919_),
    .A2(_09925_),
    .A3(_09936_),
    .B1(_09918_),
    .X(_09938_));
 o21ai_1 _14713_ (.A1(_09914_),
    .A2(_09938_),
    .B1(_09915_),
    .Y(_09939_));
 nand2b_1 _14714_ (.A_N(_09939_),
    .B(_09911_),
    .Y(_09940_));
 o21ai_1 _14715_ (.A1(net484),
    .A2(_09910_),
    .B1(_09940_),
    .Y(_09941_));
 or2_1 _14716_ (.A(_09907_),
    .B(_09908_),
    .X(_09942_));
 o21ba_1 _14717_ (.A1(_09908_),
    .A2(_09941_),
    .B1_N(_09907_),
    .X(_09943_));
 or2_1 _14718_ (.A(_09905_),
    .B(_09943_),
    .X(_09944_));
 and2_1 _14719_ (.A(net478),
    .B(_09876_),
    .X(_09945_));
 nor2_1 _14720_ (.A(_09902_),
    .B(_09945_),
    .Y(_09946_));
 and2_1 _14721_ (.A(net476),
    .B(_09904_),
    .X(_09947_));
 nand2_1 _14722_ (.A(net476),
    .B(_09904_),
    .Y(_09948_));
 a31o_1 _14723_ (.A1(_09944_),
    .A2(_09946_),
    .A3(_09948_),
    .B1(_09877_),
    .X(_09949_));
 xnor2_1 _14724_ (.A(_09278_),
    .B(_09726_),
    .Y(_09950_));
 nor2_1 _14725_ (.A(net517),
    .B(net477),
    .Y(_09951_));
 nor2_1 _14726_ (.A(net516),
    .B(_09757_),
    .Y(_09952_));
 nor2_1 _14727_ (.A(_09951_),
    .B(_09952_),
    .Y(_09953_));
 nor2_1 _14728_ (.A(net507),
    .B(net485),
    .Y(_09954_));
 nor2_1 _14729_ (.A(net503),
    .B(_09763_),
    .Y(_09955_));
 nor2_1 _14730_ (.A(_09954_),
    .B(_09955_),
    .Y(_09956_));
 nor2_1 _14731_ (.A(net497),
    .B(_09769_),
    .Y(_09957_));
 nor2_1 _14732_ (.A(_09269_),
    .B(_09770_),
    .Y(_09958_));
 nor2_1 _14733_ (.A(_09957_),
    .B(_09958_),
    .Y(_09959_));
 nor2_1 _14734_ (.A(net502),
    .B(net483),
    .Y(_09960_));
 and2_1 _14735_ (.A(net502),
    .B(net483),
    .X(_09961_));
 or2_1 _14736_ (.A(_09960_),
    .B(_09961_),
    .X(_09962_));
 nand2_1 _14737_ (.A(net509),
    .B(_09785_),
    .Y(_09963_));
 xnor2_1 _14738_ (.A(_09264_),
    .B(_09785_),
    .Y(_09964_));
 and3_1 _14739_ (.A(net523),
    .B(net489),
    .C(_09791_),
    .X(_09965_));
 a21o_1 _14740_ (.A1(net490),
    .A2(_09791_),
    .B1(net523),
    .X(_09966_));
 nand2b_1 _14741_ (.A_N(_09965_),
    .B(_09966_),
    .Y(_09967_));
 a21o_1 _14742_ (.A1(net487),
    .A2(net492),
    .B1(net512),
    .X(_09968_));
 and3b_1 _14743_ (.A_N(_09965_),
    .B(_09966_),
    .C(_09968_),
    .X(_09969_));
 o21ai_1 _14744_ (.A1(_09965_),
    .A2(_09969_),
    .B1(_09964_),
    .Y(_09970_));
 a21oi_1 _14745_ (.A1(_09963_),
    .A2(_09970_),
    .B1(_09962_),
    .Y(_09971_));
 o21a_1 _14746_ (.A1(_09960_),
    .A2(_09971_),
    .B1(_09959_),
    .X(_09972_));
 o21a_1 _14747_ (.A1(_09957_),
    .A2(_09972_),
    .B1(_09956_),
    .X(_09973_));
 o21a_1 _14748_ (.A1(_09954_),
    .A2(_09973_),
    .B1(_09953_),
    .X(_09974_));
 o21ai_1 _14749_ (.A1(_09951_),
    .A2(_09974_),
    .B1(_09950_),
    .Y(_09975_));
 o21ai_1 _14750_ (.A1(net521),
    .A2(net478),
    .B1(_09975_),
    .Y(_09976_));
 or2_1 _14751_ (.A(net520),
    .B(net485),
    .X(_09977_));
 inv_2 _14752_ (.A(_09977_),
    .Y(_09978_));
 nand2_1 _14753_ (.A(net520),
    .B(net485),
    .Y(_09979_));
 nand2_1 _14754_ (.A(_09977_),
    .B(_09979_),
    .Y(_09980_));
 nor2_1 _14755_ (.A(net519),
    .B(net484),
    .Y(_09981_));
 nand2_1 _14756_ (.A(net519),
    .B(net484),
    .Y(_09982_));
 nand2b_1 _14757_ (.A_N(_09981_),
    .B(_09982_),
    .Y(_09983_));
 nand2_1 _14758_ (.A(net504),
    .B(net482),
    .Y(_09984_));
 nor2_1 _14759_ (.A(net504),
    .B(net482),
    .Y(_09985_));
 inv_2 _14760_ (.A(_09985_),
    .Y(_09986_));
 nor2_1 _14761_ (.A(net496),
    .B(net481),
    .Y(_09987_));
 nand2_1 _14762_ (.A(net498),
    .B(net481),
    .Y(_09988_));
 nand2b_1 _14763_ (.A_N(_09987_),
    .B(_09988_),
    .Y(_09989_));
 nor2_1 _14764_ (.A(net501),
    .B(net479),
    .Y(_09990_));
 nand2_1 _14765_ (.A(net501),
    .B(net479),
    .Y(_09991_));
 a211o_1 _14766_ (.A1(_09806_),
    .A2(_09807_),
    .B1(_09990_),
    .C1(_09800_),
    .X(_09992_));
 nand2_1 _14767_ (.A(_09991_),
    .B(_09992_),
    .Y(_09993_));
 a31o_1 _14768_ (.A1(_09988_),
    .A2(_09991_),
    .A3(_09992_),
    .B1(_09987_),
    .X(_09994_));
 o21ai_1 _14769_ (.A1(_09985_),
    .A2(_09994_),
    .B1(_09984_),
    .Y(_09995_));
 nor2_1 _14770_ (.A(_09983_),
    .B(_09995_),
    .Y(_09996_));
 o31a_1 _14771_ (.A1(_09980_),
    .A2(_09981_),
    .A3(_09996_),
    .B1(net478),
    .X(_09997_));
 o21ai_1 _14772_ (.A1(_09981_),
    .A2(_09996_),
    .B1(_09980_),
    .Y(_09998_));
 and2_1 _14773_ (.A(_09983_),
    .B(_09995_),
    .X(_09999_));
 o311a_1 _14774_ (.A1(net520),
    .A2(_09996_),
    .A3(_09999_),
    .B1(_09998_),
    .C1(_09997_),
    .X(_10000_));
 nand2_1 _14775_ (.A(_09984_),
    .B(_09986_),
    .Y(_10001_));
 xor2_1 _14776_ (.A(_09994_),
    .B(_10001_),
    .X(_10002_));
 xnor2_1 _14777_ (.A(_09989_),
    .B(_09993_),
    .Y(_10003_));
 and2_1 _14778_ (.A(_09264_),
    .B(_09930_),
    .X(_10004_));
 a221oi_1 _14779_ (.A1(net522),
    .A2(net509),
    .B1(_09803_),
    .B2(_09804_),
    .C1(net513),
    .Y(_10005_));
 o31a_1 _14780_ (.A1(_09805_),
    .A2(_10004_),
    .A3(_10005_),
    .B1(net501),
    .X(_10006_));
 or4_1 _14781_ (.A(net501),
    .B(_09805_),
    .C(_10004_),
    .D(_10005_),
    .X(_10007_));
 xnor2_1 _14782_ (.A(_09806_),
    .B(_09808_),
    .Y(_10008_));
 o21ai_1 _14783_ (.A1(_10006_),
    .A2(_10008_),
    .B1(_10007_),
    .Y(_10009_));
 nand2_1 _14784_ (.A(net499),
    .B(_10009_),
    .Y(_10010_));
 nor2_1 _14785_ (.A(net499),
    .B(_10009_),
    .Y(_10011_));
 and2b_1 _14786_ (.A_N(_09990_),
    .B(_09991_),
    .X(_10012_));
 xnor2_1 _14787_ (.A(_09809_),
    .B(_10012_),
    .Y(_10013_));
 a221o_1 _14788_ (.A1(net507),
    .A2(_10003_),
    .B1(_10010_),
    .B2(_10013_),
    .C1(_10011_),
    .X(_10014_));
 o221a_1 _14789_ (.A1(net517),
    .A2(_10002_),
    .B1(_10003_),
    .B2(net506),
    .C1(_10014_),
    .X(_10015_));
 a211o_1 _14790_ (.A1(net517),
    .A2(_10002_),
    .B1(_10015_),
    .C1(_09854_),
    .X(_10016_));
 o21ai_1 _14791_ (.A1(_09978_),
    .A2(_09981_),
    .B1(_09979_),
    .Y(_10017_));
 o31a_1 _14792_ (.A1(_09980_),
    .A2(_09983_),
    .A3(_09995_),
    .B1(_10017_),
    .X(_10018_));
 xnor2_1 _14793_ (.A(_09757_),
    .B(_10018_),
    .Y(_10019_));
 nand2_1 _14794_ (.A(net505),
    .B(net484),
    .Y(_10020_));
 inv_2 _14795_ (.A(_10020_),
    .Y(_10021_));
 nor2_1 _14796_ (.A(net504),
    .B(net484),
    .Y(_10022_));
 nor2_1 _14797_ (.A(net496),
    .B(net482),
    .Y(_10023_));
 nand2_1 _14798_ (.A(net496),
    .B(net482),
    .Y(_10024_));
 nand2b_1 _14799_ (.A_N(_10023_),
    .B(_10024_),
    .Y(_10025_));
 nand2_1 _14800_ (.A(net510),
    .B(_09785_),
    .Y(_10026_));
 nand2_1 _14801_ (.A(net501),
    .B(net481),
    .Y(_10027_));
 a21oi_1 _14802_ (.A1(net487),
    .A2(net492),
    .B1(net522),
    .Y(_10028_));
 a21o_1 _14803_ (.A1(net488),
    .A2(net492),
    .B1(net522),
    .X(_10029_));
 and3_1 _14804_ (.A(net522),
    .B(net488),
    .C(net492),
    .X(_10030_));
 a21o_1 _14805_ (.A1(_07149_),
    .A2(net487),
    .B1(net512),
    .X(_10031_));
 nor2_1 _14806_ (.A(_10028_),
    .B(_10030_),
    .Y(_10032_));
 a21o_1 _14807_ (.A1(_10029_),
    .A2(_10031_),
    .B1(_10030_),
    .X(_10033_));
 xnor2_1 _14808_ (.A(net509),
    .B(net480),
    .Y(_10034_));
 a32o_1 _14809_ (.A1(net509),
    .A2(net488),
    .A3(_09791_),
    .B1(_10033_),
    .B2(_10034_),
    .X(_10035_));
 nand2b_1 _14810_ (.A_N(_10035_),
    .B(_10026_),
    .Y(_10036_));
 and2_1 _14811_ (.A(_10027_),
    .B(_10036_),
    .X(_10037_));
 a31o_1 _14812_ (.A1(_10024_),
    .A2(_10027_),
    .A3(_10036_),
    .B1(_10023_),
    .X(_10038_));
 a21oi_1 _14813_ (.A1(_10020_),
    .A2(_10038_),
    .B1(_10022_),
    .Y(_10039_));
 or2_1 _14814_ (.A(net521),
    .B(net476),
    .X(_10040_));
 inv_2 _14815_ (.A(_10040_),
    .Y(_10041_));
 nor2_1 _14816_ (.A(_09278_),
    .B(_09757_),
    .Y(_10042_));
 xnor2_1 _14817_ (.A(net517),
    .B(net485),
    .Y(_10043_));
 or4_1 _14818_ (.A(_10039_),
    .B(_10041_),
    .C(_10042_),
    .D(_10043_),
    .X(_10044_));
 o311a_1 _14819_ (.A1(net518),
    .A2(net485),
    .A3(_10042_),
    .B1(_10040_),
    .C1(net478),
    .X(_10045_));
 nand2_1 _14820_ (.A(_10044_),
    .B(_10045_),
    .Y(_10046_));
 nand2b_1 _14821_ (.A_N(_09800_),
    .B(_09803_),
    .Y(_10047_));
 a31o_1 _14822_ (.A1(net512),
    .A2(_09804_),
    .A3(_09977_),
    .B1(_10047_),
    .X(_10048_));
 a311o_1 _14823_ (.A1(_09807_),
    .A2(_09991_),
    .A3(_10048_),
    .B1(_09987_),
    .C1(_09990_),
    .X(_10049_));
 a311o_1 _14824_ (.A1(_09984_),
    .A2(_09988_),
    .A3(_10049_),
    .B1(_09985_),
    .C1(_09981_),
    .X(_10050_));
 or3_1 _14825_ (.A(_09727_),
    .B(_09757_),
    .C(_09978_),
    .X(_10051_));
 a31oi_1 _14826_ (.A1(_09979_),
    .A2(_09982_),
    .A3(_10050_),
    .B1(_10051_),
    .Y(_10052_));
 a311o_1 _14827_ (.A1(_10000_),
    .A2(_10016_),
    .A3(_10019_),
    .B1(_10046_),
    .C1(_10052_),
    .X(_10053_));
 nand2_1 _14828_ (.A(net476),
    .B(_09876_),
    .Y(_10054_));
 inv_2 _14829_ (.A(_10054_),
    .Y(_10055_));
 nor2_1 _14830_ (.A(net485),
    .B(_09880_),
    .Y(_10056_));
 nand2_1 _14831_ (.A(net485),
    .B(_09880_),
    .Y(_10057_));
 and2b_1 _14832_ (.A_N(_10056_),
    .B(_10057_),
    .X(_10058_));
 and3_1 _14833_ (.A(net490),
    .B(_09768_),
    .C(_09884_),
    .X(_10059_));
 nor2_1 _14834_ (.A(_09770_),
    .B(_09884_),
    .Y(_10060_));
 nor2_1 _14835_ (.A(_10059_),
    .B(_10060_),
    .Y(_10061_));
 nor2_1 _14836_ (.A(net482),
    .B(_09885_),
    .Y(_10062_));
 and2_1 _14837_ (.A(net482),
    .B(_09885_),
    .X(_10063_));
 or2_1 _14838_ (.A(_10062_),
    .B(_10063_),
    .X(_10064_));
 inv_2 _14839_ (.A(_10064_),
    .Y(_10065_));
 or2_1 _14840_ (.A(net481),
    .B(_09889_),
    .X(_10066_));
 nand2_1 _14841_ (.A(net481),
    .B(_09889_),
    .Y(_10067_));
 nand2_1 _14842_ (.A(_10066_),
    .B(_10067_),
    .Y(_10068_));
 nor2_1 _14843_ (.A(net479),
    .B(_09894_),
    .Y(_10069_));
 nand2_1 _14844_ (.A(net479),
    .B(_09894_),
    .Y(_10070_));
 nand2b_1 _14845_ (.A_N(_10069_),
    .B(_10070_),
    .Y(_10071_));
 and3_1 _14846_ (.A(net488),
    .B(net492),
    .C(_09927_),
    .X(_10072_));
 a21o_1 _14847_ (.A1(net488),
    .A2(_09798_),
    .B1(_09927_),
    .X(_10073_));
 and2b_1 _14848_ (.A_N(_10072_),
    .B(_10073_),
    .X(_10074_));
 a31o_1 _14849_ (.A1(_09804_),
    .A2(_09930_),
    .A3(_10073_),
    .B1(_10072_),
    .X(_10075_));
 a21o_1 _14850_ (.A1(_10070_),
    .A2(_10075_),
    .B1(_10069_),
    .X(_10076_));
 a21bo_1 _14851_ (.A1(_10067_),
    .A2(_10076_),
    .B1_N(_10066_),
    .X(_10077_));
 a21o_1 _14852_ (.A1(_10065_),
    .A2(_10077_),
    .B1(_10062_),
    .X(_10078_));
 a21o_1 _14853_ (.A1(_10061_),
    .A2(_10078_),
    .B1(_10059_),
    .X(_10079_));
 a21o_1 _14854_ (.A1(_10057_),
    .A2(_10079_),
    .B1(_10056_),
    .X(_10080_));
 o21ai_1 _14855_ (.A1(net476),
    .A2(_09876_),
    .B1(net478),
    .Y(_10081_));
 a21oi_1 _14856_ (.A1(_10054_),
    .A2(_10080_),
    .B1(_10081_),
    .Y(_10082_));
 xnor2_1 _14857_ (.A(_10025_),
    .B(_10037_),
    .Y(_10083_));
 nand2_1 _14858_ (.A(_10026_),
    .B(_10027_),
    .Y(_10084_));
 xor2_1 _14859_ (.A(_10035_),
    .B(_10084_),
    .X(_10085_));
 xnor2_1 _14860_ (.A(_10033_),
    .B(_10034_),
    .Y(_10086_));
 o21ai_1 _14861_ (.A1(_07149_),
    .A2(_09753_),
    .B1(_10031_),
    .Y(_10087_));
 a21oi_1 _14862_ (.A1(net508),
    .A2(_10087_),
    .B1(net511),
    .Y(_10088_));
 nand2_1 _14863_ (.A(_09271_),
    .B(_10087_),
    .Y(_10089_));
 xnor2_1 _14864_ (.A(_10031_),
    .B(_10032_),
    .Y(_10090_));
 a221o_1 _14865_ (.A1(net496),
    .A2(_10086_),
    .B1(_10089_),
    .B2(_10090_),
    .C1(_10088_),
    .X(_10091_));
 o221a_1 _14866_ (.A1(net505),
    .A2(_10085_),
    .B1(_10086_),
    .B2(net496),
    .C1(_10091_),
    .X(_10092_));
 a21oi_1 _14867_ (.A1(net505),
    .A2(_10085_),
    .B1(_10092_),
    .Y(_10093_));
 a21o_1 _14868_ (.A1(net515),
    .A2(_10083_),
    .B1(_10093_),
    .X(_10094_));
 o211a_1 _14869_ (.A1(net515),
    .A2(_10083_),
    .B1(_10094_),
    .C1(_09855_),
    .X(_10095_));
 o22a_1 _14870_ (.A1(net515),
    .A2(_09763_),
    .B1(_10041_),
    .B2(_10042_),
    .X(_10096_));
 or2_1 _14871_ (.A(_10021_),
    .B(_10022_),
    .X(_10097_));
 xnor2_1 _14872_ (.A(_10038_),
    .B(_10097_),
    .Y(_10098_));
 a221o_1 _14873_ (.A1(_10054_),
    .A2(_10080_),
    .B1(_10098_),
    .B2(_09278_),
    .C1(_10081_),
    .X(_10099_));
 or4b_1 _14874_ (.A(_10095_),
    .B(_10099_),
    .C(_10096_),
    .D_N(_10046_),
    .X(_10100_));
 a221o_1 _14875_ (.A1(net506),
    .A2(_09786_),
    .B1(net479),
    .B2(_09847_),
    .C1(_09849_),
    .X(_10101_));
 o221a_1 _14876_ (.A1(net517),
    .A2(net483),
    .B1(_09786_),
    .B2(net507),
    .C1(_10101_),
    .X(_10102_));
 a211o_1 _14877_ (.A1(net517),
    .A2(net483),
    .B1(_09854_),
    .C1(_10102_),
    .X(_10103_));
 o211a_1 _14878_ (.A1(net521),
    .A2(_09769_),
    .B1(_10052_),
    .C1(_10103_),
    .X(_10104_));
 inv_2 _14879_ (.A(_10104_),
    .Y(_10105_));
 xnor2_1 _14880_ (.A(_10058_),
    .B(_10079_),
    .Y(_10106_));
 xnor2_1 _14881_ (.A(_10061_),
    .B(_10078_),
    .Y(_10107_));
 xnor2_1 _14882_ (.A(_10065_),
    .B(_10077_),
    .Y(_10108_));
 xor2_1 _14883_ (.A(_10068_),
    .B(_10076_),
    .X(_10109_));
 xnor2_1 _14884_ (.A(_10071_),
    .B(_10075_),
    .Y(_10110_));
 o211a_1 _14885_ (.A1(net512),
    .A2(_09921_),
    .B1(_09804_),
    .C1(_09803_),
    .X(_10111_));
 or2_1 _14886_ (.A(_10004_),
    .B(_10111_),
    .X(_10112_));
 nor2_1 _14887_ (.A(net502),
    .B(_10112_),
    .Y(_10113_));
 nand2_1 _14888_ (.A(net502),
    .B(_10112_),
    .Y(_10114_));
 xnor2_1 _14889_ (.A(_09931_),
    .B(_10074_),
    .Y(_10115_));
 a221o_1 _14890_ (.A1(net500),
    .A2(_10110_),
    .B1(_10114_),
    .B2(_10115_),
    .C1(_10113_),
    .X(_10116_));
 o2bb2a_1 _14891_ (.A1_N(net505),
    .A2_N(_10109_),
    .B1(_10110_),
    .B2(net500),
    .X(_10117_));
 nand2_1 _14892_ (.A(_10116_),
    .B(_10117_),
    .Y(_10118_));
 o221a_1 _14893_ (.A1(net519),
    .A2(_10108_),
    .B1(_10109_),
    .B2(net504),
    .C1(_10118_),
    .X(_10119_));
 a211o_1 _14894_ (.A1(net519),
    .A2(_10108_),
    .B1(_10119_),
    .C1(_09854_),
    .X(_10120_));
 o221a_1 _14895_ (.A1(net478),
    .A2(_10055_),
    .B1(_10107_),
    .B2(net520),
    .C1(_10106_),
    .X(_10121_));
 nand2_1 _14896_ (.A(_10080_),
    .B(_10081_),
    .Y(_10122_));
 a31o_1 _14897_ (.A1(_10120_),
    .A2(_10121_),
    .A3(_10122_),
    .B1(_10082_),
    .X(_10123_));
 a41oi_1 _14898_ (.A1(_10053_),
    .A2(_10100_),
    .A3(_10105_),
    .A4(_10123_),
    .B1(_09976_),
    .Y(_10124_));
 nor2_1 _14899_ (.A(_09686_),
    .B(_09763_),
    .Y(_10125_));
 nand2_1 _14900_ (.A(_09686_),
    .B(_09763_),
    .Y(_10126_));
 and3_1 _14901_ (.A(_09688_),
    .B(net490),
    .C(_09768_),
    .X(_10127_));
 nor2_1 _14902_ (.A(_09688_),
    .B(_09770_),
    .Y(_10128_));
 nor2_1 _14903_ (.A(_10127_),
    .B(_10128_),
    .Y(_10129_));
 and3_1 _14904_ (.A(_09691_),
    .B(net490),
    .C(_09776_),
    .X(_10130_));
 a21o_1 _14905_ (.A1(net490),
    .A2(_09776_),
    .B1(_09691_),
    .X(_10131_));
 nor2_1 _14906_ (.A(_09695_),
    .B(net481),
    .Y(_10132_));
 nor2_1 _14907_ (.A(_09694_),
    .B(_09785_),
    .Y(_10133_));
 nor2_1 _14908_ (.A(_10132_),
    .B(_10133_),
    .Y(_10134_));
 nor2_1 _14909_ (.A(_09699_),
    .B(net480),
    .Y(_10135_));
 nand2_1 _14910_ (.A(_09699_),
    .B(net480),
    .Y(_10136_));
 and3_1 _14911_ (.A(_09705_),
    .B(net489),
    .C(net492),
    .X(_10137_));
 xnor2_1 _14912_ (.A(_09704_),
    .B(_09799_),
    .Y(_10138_));
 a21o_1 _14913_ (.A1(_09806_),
    .A2(_10138_),
    .B1(_10137_),
    .X(_10139_));
 a211o_1 _14914_ (.A1(_09806_),
    .A2(_10138_),
    .B1(_10137_),
    .C1(_10135_),
    .X(_10140_));
 nand2_1 _14915_ (.A(_10136_),
    .B(_10140_),
    .Y(_10141_));
 a31o_1 _14916_ (.A1(_10134_),
    .A2(_10136_),
    .A3(_10140_),
    .B1(_10132_),
    .X(_10142_));
 o21a_1 _14917_ (.A1(_10130_),
    .A2(_10142_),
    .B1(_10131_),
    .X(_10143_));
 o211a_1 _14918_ (.A1(_10130_),
    .A2(_10142_),
    .B1(_10131_),
    .C1(_10129_),
    .X(_10144_));
 a211o_1 _14919_ (.A1(_09686_),
    .A2(_09763_),
    .B1(_10127_),
    .C1(_10144_),
    .X(_10145_));
 nand2b_1 _14920_ (.A_N(_10125_),
    .B(_10145_),
    .Y(_10146_));
 nand2_1 _14921_ (.A(_09722_),
    .B(_09757_),
    .Y(_10147_));
 nand2b_1 _14922_ (.A_N(_10130_),
    .B(_10131_),
    .Y(_10148_));
 nand2b_1 _14923_ (.A_N(_10135_),
    .B(_10136_),
    .Y(_10149_));
 nand2b_1 _14924_ (.A_N(_10125_),
    .B(_10126_),
    .Y(_10150_));
 nand2_1 _14925_ (.A(_10146_),
    .B(_10147_),
    .Y(_10151_));
 or2_1 _14926_ (.A(_09722_),
    .B(_09757_),
    .X(_10152_));
 nand2_1 _14927_ (.A(_09278_),
    .B(_09720_),
    .Y(_10153_));
 a21oi_1 _14928_ (.A1(net478),
    .A2(_10153_),
    .B1(_09877_),
    .Y(_10154_));
 and3_1 _14929_ (.A(_10151_),
    .B(_10152_),
    .C(_10154_),
    .X(_10155_));
 nor2_1 _14930_ (.A(_09877_),
    .B(_10155_),
    .Y(_10156_));
 or3_1 _14931_ (.A(_09950_),
    .B(_09951_),
    .C(_09974_),
    .X(_10157_));
 or3_1 _14932_ (.A(_09953_),
    .B(_09954_),
    .C(_09973_),
    .X(_10158_));
 and2b_1 _14933_ (.A_N(_09974_),
    .B(_10158_),
    .X(_10159_));
 nor3_1 _14934_ (.A(_09956_),
    .B(_09957_),
    .C(_09972_),
    .Y(_10160_));
 nor2_1 _14935_ (.A(_09973_),
    .B(_10160_),
    .Y(_10161_));
 and3_1 _14936_ (.A(_09962_),
    .B(_09963_),
    .C(_09970_),
    .X(_10162_));
 nor2_1 _14937_ (.A(_09971_),
    .B(_10162_),
    .Y(_10163_));
 or3_1 _14938_ (.A(_09964_),
    .B(_09965_),
    .C(_09969_),
    .X(_10164_));
 nand2_1 _14939_ (.A(_09970_),
    .B(_10164_),
    .Y(_10165_));
 xor2_1 _14940_ (.A(_09967_),
    .B(_09968_),
    .X(_10166_));
 a21bo_1 _14941_ (.A1(_09271_),
    .A2(_09802_),
    .B1_N(_09968_),
    .X(_10167_));
 a21oi_1 _14942_ (.A1(net512),
    .A2(_09799_),
    .B1(_10167_),
    .Y(_10168_));
 a211o_1 _14943_ (.A1(net497),
    .A2(_10166_),
    .B1(_10168_),
    .C1(_09844_),
    .X(_10169_));
 o221ai_1 _14944_ (.A1(net506),
    .A2(_10165_),
    .B1(_10166_),
    .B2(net497),
    .C1(_10169_),
    .Y(_10170_));
 o2bb2a_1 _14945_ (.A1_N(net506),
    .A2_N(_10165_),
    .B1(net515),
    .B2(_10163_),
    .X(_10171_));
 a22o_1 _14946_ (.A1(net515),
    .A2(_10163_),
    .B1(_10170_),
    .B2(_10171_),
    .X(_10172_));
 or3_1 _14947_ (.A(_09959_),
    .B(_09960_),
    .C(_09971_),
    .X(_10173_));
 nor2_1 _14948_ (.A(net520),
    .B(_09972_),
    .Y(_10174_));
 a22o_1 _14949_ (.A1(_09855_),
    .A2(_10172_),
    .B1(_10173_),
    .B2(_10174_),
    .X(_10175_));
 a2111oi_1 _14950_ (.A1(_09975_),
    .A2(_10157_),
    .B1(_10159_),
    .C1(_10161_),
    .D1(_10175_),
    .Y(_10176_));
 or2_1 _14951_ (.A(_09877_),
    .B(_09945_),
    .X(_10177_));
 nand2_1 _14952_ (.A(net476),
    .B(_09880_),
    .Y(_10178_));
 or2_1 _14953_ (.A(net476),
    .B(_09880_),
    .X(_10179_));
 xnor2_1 _14954_ (.A(net485),
    .B(_09884_),
    .Y(_10180_));
 nor2_1 _14955_ (.A(net484),
    .B(_09885_),
    .Y(_10181_));
 nand2_1 _14956_ (.A(net484),
    .B(_09885_),
    .Y(_10182_));
 nor2_1 _14957_ (.A(net482),
    .B(_09889_),
    .Y(_10183_));
 and2_1 _14958_ (.A(net482),
    .B(_09889_),
    .X(_10184_));
 nor2_1 _14959_ (.A(_10183_),
    .B(_10184_),
    .Y(_10185_));
 nor2_1 _14960_ (.A(net481),
    .B(_09894_),
    .Y(_10186_));
 nand2_1 _14961_ (.A(net481),
    .B(_09894_),
    .Y(_10187_));
 and3_1 _14962_ (.A(net487),
    .B(_09791_),
    .C(_09927_),
    .X(_10188_));
 a21oi_1 _14963_ (.A1(net487),
    .A2(_09791_),
    .B1(_09927_),
    .Y(_10189_));
 nor2_1 _14964_ (.A(_10188_),
    .B(_10189_),
    .Y(_10190_));
 nand2_1 _14965_ (.A(_09229_),
    .B(net514),
    .Y(_10191_));
 and2b_1 _14966_ (.A_N(_09926_),
    .B(_10191_),
    .X(_10192_));
 nand2b_1 _14967_ (.A_N(_09926_),
    .B(_10191_),
    .Y(_10193_));
 and3_1 _14968_ (.A(net487),
    .B(net492),
    .C(_10193_),
    .X(_10194_));
 a21o_1 _14969_ (.A1(net487),
    .A2(net492),
    .B1(_10193_),
    .X(_10195_));
 nand2_1 _14970_ (.A(_10031_),
    .B(_10195_),
    .Y(_10196_));
 a21o_1 _14971_ (.A1(_10031_),
    .A2(_10195_),
    .B1(_10194_),
    .X(_10197_));
 a21oi_1 _14972_ (.A1(_10190_),
    .A2(_10197_),
    .B1(_10188_),
    .Y(_10198_));
 a211o_1 _14973_ (.A1(_10190_),
    .A2(_10197_),
    .B1(_10186_),
    .C1(_10188_),
    .X(_10199_));
 nand2_1 _14974_ (.A(_10187_),
    .B(_10199_),
    .Y(_10200_));
 a31o_1 _14975_ (.A1(_10185_),
    .A2(_10187_),
    .A3(_10199_),
    .B1(_10183_),
    .X(_10201_));
 o21a_1 _14976_ (.A1(_10181_),
    .A2(_10201_),
    .B1(_10182_),
    .X(_10202_));
 o211a_1 _14977_ (.A1(_10181_),
    .A2(_10201_),
    .B1(_10182_),
    .C1(_10180_),
    .X(_10203_));
 a21o_1 _14978_ (.A1(_09763_),
    .A2(_09884_),
    .B1(_10203_),
    .X(_10204_));
 nand2_1 _14979_ (.A(_10178_),
    .B(_10204_),
    .Y(_10205_));
 a21oi_1 _14980_ (.A1(_10179_),
    .A2(_10205_),
    .B1(_10177_),
    .Y(_10206_));
 nand2_1 _14981_ (.A(_10178_),
    .B(_10179_),
    .Y(_10207_));
 nand2b_1 _14982_ (.A_N(_10186_),
    .B(_10187_),
    .Y(_10208_));
 and2b_1 _14983_ (.A_N(_10181_),
    .B(_10182_),
    .X(_10209_));
 or2_1 _14984_ (.A(_09877_),
    .B(_10206_),
    .X(_10210_));
 a31o_1 _14985_ (.A1(_10145_),
    .A2(_10147_),
    .A3(_10152_),
    .B1(_10125_),
    .X(_10211_));
 xor2_1 _14986_ (.A(_10142_),
    .B(_10148_),
    .X(_10212_));
 xor2_1 _14987_ (.A(_10134_),
    .B(_10141_),
    .X(_10213_));
 xnor2_1 _14988_ (.A(_10139_),
    .B(_10149_),
    .Y(_10214_));
 xnor2_1 _14989_ (.A(_09806_),
    .B(_10138_),
    .Y(_10215_));
 o2bb2a_1 _14990_ (.A1_N(net499),
    .A2_N(_10214_),
    .B1(_10215_),
    .B2(_10006_),
    .X(_10216_));
 nor2_1 _14991_ (.A(net499),
    .B(_10214_),
    .Y(_10217_));
 a221o_1 _14992_ (.A1(net506),
    .A2(_10213_),
    .B1(_10216_),
    .B2(_10007_),
    .C1(_10217_),
    .X(_10218_));
 o221a_1 _14993_ (.A1(net517),
    .A2(_10212_),
    .B1(_10213_),
    .B2(net507),
    .C1(_10218_),
    .X(_10219_));
 a211o_1 _14994_ (.A1(net517),
    .A2(_10212_),
    .B1(_10219_),
    .C1(_09854_),
    .X(_10220_));
 nand2_1 _14995_ (.A(_10125_),
    .B(_10147_),
    .Y(_10221_));
 o21ai_1 _14996_ (.A1(_10127_),
    .A2(_10144_),
    .B1(_10150_),
    .Y(_10222_));
 nor2_1 _14997_ (.A(_10129_),
    .B(_10143_),
    .Y(_10223_));
 o311a_1 _14998_ (.A1(net521),
    .A2(_10144_),
    .A3(_10223_),
    .B1(_10222_),
    .C1(_10154_),
    .X(_10224_));
 and4_1 _14999_ (.A(_10211_),
    .B(_10220_),
    .C(_10221_),
    .D(_10224_),
    .X(_10225_));
 nor2_1 _15000_ (.A(_10210_),
    .B(_10225_),
    .Y(_10226_));
 o41ai_1 _15001_ (.A1(_09877_),
    .A2(_10124_),
    .A3(_10155_),
    .A4(net474),
    .B1(_10226_),
    .Y(_10227_));
 and3_1 _15002_ (.A(_10177_),
    .B(_10179_),
    .C(_10205_),
    .X(_10228_));
 o21ai_1 _15003_ (.A1(_10201_),
    .A2(_10209_),
    .B1(_09278_),
    .Y(_10229_));
 a21o_1 _15004_ (.A1(_10201_),
    .A2(_10209_),
    .B1(_10229_),
    .X(_10230_));
 xnor2_1 _15005_ (.A(_10185_),
    .B(_10200_),
    .Y(_10231_));
 xnor2_1 _15006_ (.A(_10198_),
    .B(_10208_),
    .Y(_10232_));
 nand2_1 _15007_ (.A(net505),
    .B(_10232_),
    .Y(_10233_));
 xnor2_1 _15008_ (.A(_10190_),
    .B(_10197_),
    .Y(_10234_));
 o32ai_1 _15009_ (.A1(_10028_),
    .A2(_10030_),
    .A3(_10031_),
    .B1(_10194_),
    .B2(_10196_),
    .Y(_10235_));
 a221o_1 _15010_ (.A1(net496),
    .A2(_10234_),
    .B1(_10235_),
    .B2(_10089_),
    .C1(_10088_),
    .X(_10236_));
 o221ai_1 _15011_ (.A1(net505),
    .A2(_10232_),
    .B1(_10234_),
    .B2(net496),
    .C1(_10236_),
    .Y(_10237_));
 a22o_1 _15012_ (.A1(net515),
    .A2(_10231_),
    .B1(_10233_),
    .B2(_10237_),
    .X(_10238_));
 o211ai_1 _15013_ (.A1(net515),
    .A2(_10231_),
    .B1(_10238_),
    .C1(_09855_),
    .Y(_10239_));
 nor2_1 _15014_ (.A(_10180_),
    .B(_10202_),
    .Y(_10240_));
 o211a_1 _15015_ (.A1(_10203_),
    .A2(_10240_),
    .B1(_10239_),
    .C1(_10230_),
    .X(_10241_));
 xor2_1 _15016_ (.A(_10204_),
    .B(_10207_),
    .X(_10242_));
 o211ai_1 _15017_ (.A1(_10206_),
    .A2(_10228_),
    .B1(_10241_),
    .C1(_10242_),
    .Y(_10243_));
 a21oi_1 _15018_ (.A1(_10227_),
    .A2(_10243_),
    .B1(_09949_),
    .Y(_10244_));
 nor2_1 _15019_ (.A(_09839_),
    .B(_09949_),
    .Y(_10245_));
 and2b_1 _15020_ (.A_N(_09947_),
    .B(_09877_),
    .X(_10246_));
 o22a_1 _15021_ (.A1(_09877_),
    .A2(_09905_),
    .B1(_09943_),
    .B2(_10246_),
    .X(_10247_));
 xnor2_1 _15022_ (.A(_09911_),
    .B(_09939_),
    .Y(_10248_));
 a221o_1 _15023_ (.A1(_09941_),
    .A2(_09942_),
    .B1(_10248_),
    .B2(_09278_),
    .C1(_09839_),
    .X(_10249_));
 and2b_1 _15024_ (.A_N(_09914_),
    .B(_09915_),
    .X(_10250_));
 xor2_1 _15025_ (.A(_09938_),
    .B(_10250_),
    .X(_10251_));
 nand2_1 _15026_ (.A(_09931_),
    .B(_09933_),
    .Y(_10252_));
 a31o_1 _15027_ (.A1(_09934_),
    .A2(_10114_),
    .A3(_10252_),
    .B1(_10113_),
    .X(_10253_));
 a21oi_1 _15028_ (.A1(_09924_),
    .A2(_09925_),
    .B1(_09935_),
    .Y(_10254_));
 and3_1 _15029_ (.A(_09924_),
    .B(_09925_),
    .C(_09935_),
    .X(_10255_));
 xnor2_1 _15030_ (.A(_09920_),
    .B(_09937_),
    .Y(_10256_));
 a211o_1 _15031_ (.A1(net500),
    .A2(_10253_),
    .B1(_10254_),
    .C1(_10255_),
    .X(_10257_));
 o2bb2a_1 _15032_ (.A1_N(net504),
    .A2_N(_10256_),
    .B1(_10253_),
    .B2(net500),
    .X(_10258_));
 a2bb2o_1 _15033_ (.A1_N(net504),
    .A2_N(_10256_),
    .B1(net515),
    .B2(_10251_),
    .X(_10259_));
 a21o_1 _15034_ (.A1(_10257_),
    .A2(_10258_),
    .B1(_10259_),
    .X(_10260_));
 o211a_1 _15035_ (.A1(net515),
    .A2(_10251_),
    .B1(_10260_),
    .C1(_09855_),
    .X(_10261_));
 or2_1 _15036_ (.A(_09941_),
    .B(_09942_),
    .X(_10262_));
 or4b_1 _15037_ (.A(_10247_),
    .B(_10249_),
    .C(_10261_),
    .D_N(_10262_),
    .X(_10263_));
 o21a_1 _15038_ (.A1(_09839_),
    .A2(_09949_),
    .B1(_10263_),
    .X(_10264_));
 o21ba_1 _15039_ (.A1(_10244_),
    .A2(_10264_),
    .B1_N(_09860_),
    .X(_10265_));
 xnor2_1 _15040_ (.A(_09814_),
    .B(_09816_),
    .Y(_10266_));
 xnor2_1 _15041_ (.A(_09782_),
    .B(_09812_),
    .Y(_10267_));
 xnor2_1 _15042_ (.A(net513),
    .B(_10013_),
    .Y(_10268_));
 xnor2_1 _15043_ (.A(_09789_),
    .B(_09811_),
    .Y(_10269_));
 a221o_1 _15044_ (.A1(_10010_),
    .A2(_10268_),
    .B1(_10269_),
    .B2(net506),
    .C1(_10011_),
    .X(_10270_));
 o221a_1 _15045_ (.A1(net517),
    .A2(_10267_),
    .B1(_10269_),
    .B2(net507),
    .C1(_10270_),
    .X(_10271_));
 a211o_1 _15046_ (.A1(net517),
    .A2(_10267_),
    .B1(_10271_),
    .C1(_09854_),
    .X(_10272_));
 xnor2_1 _15047_ (.A(_09775_),
    .B(_09813_),
    .Y(_10273_));
 o32a_1 _15048_ (.A1(_09726_),
    .A2(_09741_),
    .A3(_09819_),
    .B1(_10273_),
    .B2(net520),
    .X(_10274_));
 nand2_1 _15049_ (.A(_10272_),
    .B(_10274_),
    .Y(_10275_));
 a211o_1 _15050_ (.A1(_09760_),
    .A2(_09817_),
    .B1(_10266_),
    .C1(_10275_),
    .X(_10276_));
 and2_1 _15051_ (.A(_09695_),
    .B(net483),
    .X(_10277_));
 o21ba_1 _15052_ (.A1(_09704_),
    .A2(net480),
    .B1_N(_10033_),
    .X(_10278_));
 a221o_1 _15053_ (.A1(_09699_),
    .A2(_09786_),
    .B1(net480),
    .B2(_09704_),
    .C1(_10278_),
    .X(_10279_));
 o221a_1 _15054_ (.A1(_09695_),
    .A2(net483),
    .B1(_09786_),
    .B2(_09699_),
    .C1(_10279_),
    .X(_10280_));
 a2bb2o_1 _15055_ (.A1_N(_10277_),
    .A2_N(_10280_),
    .B1(_09691_),
    .B2(_09770_),
    .X(_10281_));
 o221a_1 _15056_ (.A1(_09688_),
    .A2(_09763_),
    .B1(_09770_),
    .B2(_09691_),
    .C1(_10281_),
    .X(_10282_));
 a221o_1 _15057_ (.A1(_09686_),
    .A2(_09757_),
    .B1(_09763_),
    .B2(_09688_),
    .C1(_10282_),
    .X(_10283_));
 or2_1 _15058_ (.A(_09686_),
    .B(_09757_),
    .X(_10284_));
 a31o_1 _15059_ (.A1(_09722_),
    .A2(_10283_),
    .A3(_10284_),
    .B1(_09727_),
    .X(_10285_));
 a31oi_1 _15060_ (.A1(_09742_),
    .A2(_09820_),
    .A3(_10276_),
    .B1(_09753_),
    .Y(_10286_));
 or3b_2 _15061_ (.A(_10265_),
    .B(_10285_),
    .C_N(_10286_),
    .X(_10287_));
 nor2_1 _15062_ (.A(_09860_),
    .B(_10285_),
    .Y(_10288_));
 or2_1 _15063_ (.A(_09860_),
    .B(_10285_),
    .X(_10289_));
 nor2_1 _15064_ (.A(_09753_),
    .B(_10288_),
    .Y(_10290_));
 or2_1 _15065_ (.A(_10046_),
    .B(_10104_),
    .X(_10291_));
 and3b_1 _15066_ (.A_N(_09976_),
    .B(_10100_),
    .C(_10291_),
    .X(_10292_));
 o21ai_1 _15067_ (.A1(net474),
    .A2(_10292_),
    .B1(_10156_),
    .Y(_10293_));
 nand2_1 _15068_ (.A(_10210_),
    .B(_10243_),
    .Y(_10294_));
 a41o_1 _15069_ (.A1(net490),
    .A2(_10245_),
    .A3(_10293_),
    .A4(_10294_),
    .B1(_10290_),
    .X(_10295_));
 inv_2 _15070_ (.A(_10295_),
    .Y(_10296_));
 and4bb_1 _15071_ (.A_N(_10265_),
    .B_N(_10285_),
    .C(_10286_),
    .D(_10295_),
    .X(_10297_));
 or4_1 _15072_ (.A(_09839_),
    .B(_09949_),
    .C(_09976_),
    .D(_10155_),
    .X(_10298_));
 nor2_1 _15073_ (.A(_10104_),
    .B(_10298_),
    .Y(_10299_));
 a31o_1 _15074_ (.A1(_10156_),
    .A2(_10176_),
    .A3(_10245_),
    .B1(_10289_),
    .X(_10300_));
 o21ai_2 _15075_ (.A1(_10299_),
    .A2(_10300_),
    .B1(net490),
    .Y(_10301_));
 xnor2_1 _15076_ (.A(_10297_),
    .B(_10301_),
    .Y(_10302_));
 o31a_1 _15077_ (.A1(_09753_),
    .A2(_10288_),
    .A3(_10297_),
    .B1(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[4] ),
    .X(_10303_));
 xnor2_1 _15078_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[2] ),
    .B(_10302_),
    .Y(_10304_));
 o211ai_1 _15079_ (.A1(_10105_),
    .A2(_10298_),
    .B1(_10288_),
    .C1(net490),
    .Y(_10305_));
 or4_1 _15080_ (.A(_10287_),
    .B(_10289_),
    .C(_10296_),
    .D(_10301_),
    .X(_10306_));
 o31ai_1 _15081_ (.A1(_10287_),
    .A2(_10296_),
    .A3(_10301_),
    .B1(_10305_),
    .Y(_10307_));
 a21oi_1 _15082_ (.A1(_10306_),
    .A2(_10307_),
    .B1(_07157_),
    .Y(_10308_));
 o211a_1 _15083_ (.A1(_10287_),
    .A2(_10301_),
    .B1(_10290_),
    .C1(_07158_),
    .X(_10309_));
 xnor2_1 _15084_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[1] ),
    .B(_10295_),
    .Y(_10310_));
 nand2_1 _15085_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[0] ),
    .B(_10310_),
    .Y(_10311_));
 or2_1 _15086_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[0] ),
    .B(_10310_),
    .X(_10312_));
 mux2_1 _15087_ (.A0(_10311_),
    .A1(_10312_),
    .S(_10287_),
    .X(_10313_));
 a311o_1 _15088_ (.A1(_07157_),
    .A2(_10306_),
    .A3(_10307_),
    .B1(_10309_),
    .C1(_10313_),
    .X(_10314_));
 or4_4 _15089_ (.A(_10303_),
    .B(_10304_),
    .C(_10308_),
    .D(_10314_),
    .X(_10315_));
 inv_2 _15090_ (.A(_10315_),
    .Y(\digitop_pav2.proc_ctrl_inst.cmdfsm.n_pass_t1_i ));
 nand2_1 _15091_ (.A(\digitop_pav2.func_reg_wr_en ),
    .B(_09571_),
    .Y(_10316_));
 and3_1 _15092_ (.A(\digitop_pav2.func_reg_wr_en ),
    .B(\digitop_pav2.memctrl_inst.state[2] ),
    .C(_09571_),
    .X(_10317_));
 o31a_1 _15093_ (.A1(\digitop_pav2.memctrl_inst.ctr[7] ),
    .A2(_09570_),
    .A3(_09572_),
    .B1(\digitop_pav2.memctrl_inst.state[4] ),
    .X(_10318_));
 or4_1 _15094_ (.A(\digitop_pav2.memctrl_inst.bit_addr[0] ),
    .B(\digitop_pav2.memctrl_inst.bit_addr[1] ),
    .C(\digitop_pav2.memctrl_inst.bit_addr[3] ),
    .D(\digitop_pav2.memctrl_inst.bit_addr[2] ),
    .X(_10319_));
 a221o_1 _15095_ (.A1(\digitop_pav2.memctrl_inst.reg_wr_ok_ff2 ),
    .A2(_10317_),
    .B1(_10319_),
    .B2(\digitop_pav2.memctrl_inst.state[1] ),
    .C1(_10318_),
    .X(_00081_));
 a31o_1 _15096_ (.A1(\digitop_pav2.memctrl_inst.nvm_rd_en_i ),
    .A2(\digitop_pav2.memctrl_inst.state[0] ),
    .A3(_07929_),
    .B1(\digitop_pav2.memctrl_inst.n_read ),
    .X(_00080_));
 and3_1 _15097_ (.A(\digitop_pav2.memctrl_inst.nvm_wr_en_i ),
    .B(\digitop_pav2.memctrl_inst.state[0] ),
    .C(_07929_),
    .X(_10320_));
 nand2_1 _15098_ (.A(\digitop_pav2.memctrl_inst.state[0] ),
    .B(_07930_),
    .Y(_10321_));
 a2bb2o_1 _15099_ (.A1_N(\digitop_pav2.memctrl_inst.nvm_rd_en_i ),
    .A2_N(_10321_),
    .B1(_10316_),
    .B2(\digitop_pav2.memctrl_inst.state[2] ),
    .X(_00079_));
 nor2_1 _15100_ (.A(_07140_),
    .B(_10319_),
    .Y(_10322_));
 a31o_1 _15101_ (.A1(\digitop_pav2.func_rr_read ),
    .A2(\digitop_pav2.memctrl_inst.state[3] ),
    .A3(_09571_),
    .B1(_10322_),
    .X(_10323_));
 a211o_1 _15102_ (.A1(_07141_),
    .A2(_10317_),
    .B1(_10323_),
    .C1(_09421_),
    .X(_00078_));
 a21oi_1 _15103_ (.A1(net1176),
    .A2(_07135_),
    .B1(_07063_),
    .Y(_10324_));
 and2_1 _15104_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[3] ),
    .B(_10324_),
    .X(_10325_));
 nand2_2 _15105_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[3] ),
    .B(_10324_),
    .Y(_10326_));
 nor2_1 _15106_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[5] ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.state[1] ),
    .Y(_10327_));
 or2_1 _15107_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[5] ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.state[1] ),
    .X(_10328_));
 a31o_1 _15108_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[10] ),
    .A2(net1014),
    .A3(_10327_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.r_invent3_o ),
    .X(_00068_));
 nand2_1 _15109_ (.A(net159),
    .B(net1014),
    .Y(_10329_));
 o21ai_1 _15110_ (.A1(_07861_),
    .A2(_07868_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.state[11] ),
    .Y(_10330_));
 a2bb2o_1 _15111_ (.A1_N(_10329_),
    .A2_N(_10330_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.state[12] ),
    .B2(_10326_),
    .X(_00067_));
 a22o_1 _15112_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[4] ),
    .A2(net1014),
    .B1(_10329_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.state[11] ),
    .X(_00066_));
 nand2_1 _15113_ (.A(net1248),
    .B(net1014),
    .Y(_10331_));
 a2bb2o_1 _15114_ (.A1_N(_07131_),
    .A2_N(_10331_),
    .B1(_10326_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.state[10] ),
    .X(_00065_));
 a41o_1 _15115_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[11] ),
    .A2(net159),
    .A3(_07860_),
    .A4(_07867_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.state[12] ),
    .X(_10332_));
 nand2_2 _15116_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[3] ),
    .B(_07135_),
    .Y(_10333_));
 and2b_1 _15117_ (.A_N(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[0] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[1] ),
    .X(_10334_));
 nand2_2 _15118_ (.A(_07134_),
    .B(_10334_),
    .Y(_10335_));
 nor2_1 _15119_ (.A(_10333_),
    .B(_10335_),
    .Y(_10336_));
 and3_1 _15120_ (.A(net1691),
    .B(_07132_),
    .C(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[6] ),
    .X(_10337_));
 and4b_1 _15121_ (.A_N(_08964_),
    .B(_10336_),
    .C(_10337_),
    .D(\digitop_pav2.invent_inst.invent_sel_pav2.state[0] ),
    .X(_10338_));
 or3_2 _15122_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[0] ),
    .B(net1177),
    .C(_07134_),
    .X(_10339_));
 nand2_1 _15123_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[3] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[4] ),
    .Y(_10340_));
 nor2_1 _15124_ (.A(_10339_),
    .B(_10340_),
    .Y(_10341_));
 or2_1 _15125_ (.A(_10339_),
    .B(_10340_),
    .X(_10342_));
 o21a_1 _15126_ (.A1(_10326_),
    .A2(_10342_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.state[9] ),
    .X(_10343_));
 a211o_1 _15127_ (.A1(net1014),
    .A2(_10332_),
    .B1(_10338_),
    .C1(_10343_),
    .X(_00077_));
 and3_1 _15128_ (.A(net1691),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[7] ),
    .C(_07133_),
    .X(_10344_));
 nor2_1 _15129_ (.A(_10337_),
    .B(_10344_),
    .Y(_10345_));
 or2_1 _15130_ (.A(_08964_),
    .B(_10345_),
    .X(_10346_));
 a41o_1 _15131_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[0] ),
    .A2(net1014),
    .A3(_10336_),
    .A4(_10346_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.r_invent2_o ),
    .X(_00076_));
 nand2_1 _15132_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[0] ),
    .B(_07860_),
    .Y(_10347_));
 or2_1 _15133_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[0] ),
    .B(_07860_),
    .X(_10348_));
 nand2_1 _15134_ (.A(_10347_),
    .B(_10348_),
    .Y(_10349_));
 and3_1 _15135_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[2] ),
    .B(net1271),
    .C(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[2] ),
    .X(_10350_));
 and3_1 _15136_ (.A(net1271),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[3] ),
    .C(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[3] ),
    .X(_10351_));
 a21oi_1 _15137_ (.A1(net1271),
    .A2(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[3] ),
    .B1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[3] ),
    .Y(_10352_));
 or2_1 _15138_ (.A(_10351_),
    .B(_10352_),
    .X(_10353_));
 and3_1 _15139_ (.A(net1271),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[4] ),
    .C(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[4] ),
    .X(_10354_));
 a21oi_1 _15140_ (.A1(net1271),
    .A2(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[4] ),
    .B1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[4] ),
    .Y(_10355_));
 or2_1 _15141_ (.A(_10354_),
    .B(_10355_),
    .X(_10356_));
 xor2_1 _15142_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[5] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[5] ),
    .X(_10357_));
 nand2_1 _15143_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[6] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[6] ),
    .Y(_10358_));
 and3_1 _15144_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[6] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[6] ),
    .C(_10357_),
    .X(_10359_));
 a21oi_1 _15145_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[5] ),
    .A2(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[5] ),
    .B1(_10359_),
    .Y(_10360_));
 o21bai_1 _15146_ (.A1(_10355_),
    .A2(_10360_),
    .B1_N(_10354_),
    .Y(_10361_));
 and2b_1 _15147_ (.A_N(_10353_),
    .B(_10361_),
    .X(_10362_));
 or2_1 _15148_ (.A(_10351_),
    .B(_10362_),
    .X(_10363_));
 nor2_1 _15149_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[2] ),
    .B(_07857_),
    .Y(_10364_));
 nor2_1 _15150_ (.A(_10350_),
    .B(_10364_),
    .Y(_10365_));
 a21o_1 _15151_ (.A1(_10363_),
    .A2(_10365_),
    .B1(_10350_),
    .X(_10366_));
 a21o_1 _15152_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[1] ),
    .A2(_07858_),
    .B1(_10366_),
    .X(_10367_));
 o21a_1 _15153_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[1] ),
    .A2(_07858_),
    .B1(_10367_),
    .X(_10368_));
 nand2b_1 _15154_ (.A_N(_10349_),
    .B(_10368_),
    .Y(_10369_));
 a21oi_1 _15155_ (.A1(_10347_),
    .A2(_10369_),
    .B1(_07138_),
    .Y(_10370_));
 a21o_1 _15156_ (.A1(_10347_),
    .A2(_10369_),
    .B1(_07138_),
    .X(_10371_));
 and3_1 _15157_ (.A(_07138_),
    .B(_10347_),
    .C(_10369_),
    .X(_10372_));
 nor2_1 _15158_ (.A(_10370_),
    .B(_10372_),
    .Y(_10373_));
 xor2_1 _15159_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[7] ),
    .B(_10373_),
    .X(_10374_));
 xnor2_2 _15160_ (.A(_10349_),
    .B(_10368_),
    .Y(_10375_));
 inv_2 _15161_ (.A(_10375_),
    .Y(_10376_));
 xnor2_1 _15162_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[1] ),
    .B(_07858_),
    .Y(_10377_));
 xnor2_1 _15163_ (.A(_10366_),
    .B(_10377_),
    .Y(_10378_));
 xnor2_1 _15164_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[5] ),
    .B(_10378_),
    .Y(_10379_));
 xnor2_1 _15165_ (.A(_10363_),
    .B(_10365_),
    .Y(_10380_));
 or2_1 _15166_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[4] ),
    .B(_10380_),
    .X(_10381_));
 xor2_1 _15167_ (.A(_10353_),
    .B(_10361_),
    .X(_10382_));
 xnor2_1 _15168_ (.A(_10356_),
    .B(_10360_),
    .Y(_10383_));
 nand2_1 _15169_ (.A(net1174),
    .B(_10383_),
    .Y(_10384_));
 and2b_1 _15170_ (.A_N(_10357_),
    .B(_10358_),
    .X(_10385_));
 or2_1 _15171_ (.A(_10359_),
    .B(_10385_),
    .X(_10386_));
 or2_1 _15172_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[6] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[6] ),
    .X(_10387_));
 nand2_1 _15173_ (.A(_10358_),
    .B(_10387_),
    .Y(_10388_));
 xnor2_1 _15174_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[0] ),
    .B(_10388_),
    .Y(_10389_));
 a21oi_1 _15175_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[1] ),
    .A2(_10386_),
    .B1(_10389_),
    .Y(_10390_));
 o221a_1 _15176_ (.A1(net1174),
    .A2(_10383_),
    .B1(_10386_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[1] ),
    .C1(_10390_),
    .X(_10391_));
 o211ai_1 _15177_ (.A1(net1173),
    .A2(_10382_),
    .B1(_10384_),
    .C1(_10391_),
    .Y(_10392_));
 a221oi_1 _15178_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[4] ),
    .A2(_10380_),
    .B1(_10382_),
    .B2(net1173),
    .C1(_10392_),
    .Y(_10393_));
 xor2_1 _15179_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[6] ),
    .B(_10375_),
    .X(_10394_));
 and2_1 _15180_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[8] ),
    .B(_10371_),
    .X(_10395_));
 o2111a_1 _15181_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[8] ),
    .A2(_10371_),
    .B1(_10379_),
    .C1(_10381_),
    .D1(_10393_),
    .X(_10396_));
 or4b_2 _15182_ (.A(_10374_),
    .B(_10394_),
    .C(_10395_),
    .D_N(_10396_),
    .X(_10397_));
 nor2_1 _15183_ (.A(_10342_),
    .B(_10397_),
    .Y(_10398_));
 o211a_1 _15184_ (.A1(_10342_),
    .A2(_10397_),
    .B1(_07128_),
    .C1(net1014),
    .X(_10399_));
 or2_1 _15185_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[0] ),
    .B(net1175),
    .X(_10400_));
 or2_2 _15186_ (.A(net1174),
    .B(net1173),
    .X(_10401_));
 nor2_2 _15187_ (.A(_10400_),
    .B(_10401_),
    .Y(_10402_));
 or2_1 _15188_ (.A(_10400_),
    .B(_10401_),
    .X(_10403_));
 or3_1 _15189_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[4] ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[5] ),
    .C(_10403_),
    .X(_10404_));
 xor2_1 _15190_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[6] ),
    .B(_10404_),
    .X(_10405_));
 o21ai_1 _15191_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[4] ),
    .A2(_10403_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[5] ),
    .Y(_10406_));
 and2_1 _15192_ (.A(_10404_),
    .B(_10406_),
    .X(_10407_));
 or2_2 _15193_ (.A(_07137_),
    .B(net1175),
    .X(_10408_));
 nand2b_2 _15194_ (.A_N(net1174),
    .B(net1173),
    .Y(_10409_));
 nor2_2 _15195_ (.A(_10408_),
    .B(_10409_),
    .Y(_10410_));
 xnor2_2 _15196_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[4] ),
    .B(_10402_),
    .Y(_10411_));
 or4bb_1 _15197_ (.A(_10407_),
    .B(_10411_),
    .C_N(_10410_),
    .D_N(_10405_),
    .X(_10412_));
 inv_2 _15198_ (.A(_10412_),
    .Y(_10413_));
 a211o_1 _15199_ (.A1(_07900_),
    .A2(_10413_),
    .B1(_10398_),
    .C1(\digitop_pav2.invent_inst.invent_sel_pav2.mask_mismatch_ff ),
    .X(_10414_));
 nand2_1 _15200_ (.A(net1014),
    .B(_10414_),
    .Y(_10415_));
 a22o_1 _15201_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[6] ),
    .A2(_10399_),
    .B1(_10415_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.state[7] ),
    .X(_00075_));
 and3_1 _15202_ (.A(net1238),
    .B(\digitop_pav2.access_inst.access_ctrl0.state[0] ),
    .C(_07395_),
    .X(_10416_));
 o211a_1 _15203_ (.A1(net1239),
    .A2(_07418_),
    .B1(_07481_),
    .C1(_10416_),
    .X(_00014_));
 nor2_1 _15204_ (.A(_07107_),
    .B(\digitop_pav2.sec_inst.sm.st[6] ),
    .Y(_10417_));
 or2_1 _15205_ (.A(_07107_),
    .B(\digitop_pav2.sec_inst.sm.st[6] ),
    .X(_10418_));
 or2_2 _15206_ (.A(net718),
    .B(net602),
    .X(_10419_));
 a211oi_2 _15207_ (.A1(net715),
    .A2(\digitop_pav2.sec_inst.ld_mem.st[2] ),
    .B1(net1033),
    .C1(_10419_),
    .Y(_10420_));
 a211o_1 _15208_ (.A1(net715),
    .A2(\digitop_pav2.sec_inst.ld_mem.st[2] ),
    .B1(net1033),
    .C1(_10419_),
    .X(_10421_));
 or4b_2 _15209_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[2] ),
    .B(_07040_),
    .C(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[0] ),
    .D_N(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[3] ),
    .X(_10422_));
 inv_2 _15210_ (.A(_10422_),
    .Y(_10423_));
 a32o_1 _15211_ (.A1(net426),
    .A2(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_2b_o ),
    .A3(_10423_),
    .B1(_10420_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[0] ),
    .X(_00043_));
 mux2_1 _15212_ (.A0(\digitop_pav2.access_inst.access_ctrl0.state[9] ),
    .A1(\digitop_pav2.access_inst.access_ctrl0.state[2] ),
    .S(_07960_),
    .X(_00032_));
 or3b_1 _15213_ (.A(net1260),
    .B(\digitop_pav2.access_inst.access_ctrl0.nvm_busy_i ),
    .C_N(\digitop_pav2.access_inst.access_ctrl0.state[10] ),
    .X(_10424_));
 or3b_1 _15214_ (.A(net1206),
    .B(_10424_),
    .C_N(_07505_),
    .X(_10425_));
 o21ai_1 _15215_ (.A1(_07091_),
    .A2(net1190),
    .B1(_10425_),
    .Y(_00033_));
 a22o_1 _15216_ (.A1(net1148),
    .A2(net1204),
    .B1(_07959_),
    .B2(\digitop_pav2.access_inst.access_ctrl0.state[18] ),
    .X(_00034_));
 nor2_4 _15217_ (.A(net1237),
    .B(net1234),
    .Y(_10426_));
 nand2_2 _15218_ (.A(net1702),
    .B(net1650),
    .Y(_10427_));
 and4_1 _15219_ (.A(\digitop_pav2.access_inst.access_check0.pc_lock_check_sync_o ),
    .B(\digitop_pav2.access_inst.access_check0.pc_lock_check_i ),
    .C(_09522_),
    .D(_10426_),
    .X(_10428_));
 and4_1 _15220_ (.A(\digitop_pav2.access_inst.access_check0.mem_sign_check_sync_o ),
    .B(net1650),
    .C(_07970_),
    .D(_07987_),
    .X(_10429_));
 and3_1 _15221_ (.A(\digitop_pav2.access_inst.access_check0.pc_lock_check_sync_o ),
    .B(net1700),
    .C(net1192),
    .X(_10430_));
 a21o_1 _15222_ (.A1(_09522_),
    .A2(_10430_),
    .B1(_09519_),
    .X(_10431_));
 and3b_1 _15223_ (.A_N(_09523_),
    .B(_10431_),
    .C(_09518_),
    .X(_10432_));
 a2111o_1 _15224_ (.A1(\digitop_pav2.access_inst.access_ctrl0.state[5] ),
    .A2(net1207),
    .B1(_10428_),
    .C1(_10429_),
    .D1(_10432_),
    .X(_10433_));
 o21bai_1 _15225_ (.A1(_08041_),
    .A2(_08469_),
    .B1_N(_10433_),
    .Y(_00035_));
 mux2_1 _15226_ (.A0(net1063),
    .A1(\digitop_pav2.access_inst.access_ctrl0.ld_key_env_finish_i ),
    .S(\digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt ),
    .X(_10434_));
 inv_2 _15227_ (.A(_10434_),
    .Y(_10435_));
 a32o_1 _15228_ (.A1(_07023_),
    .A2(net1144),
    .A3(net1190),
    .B1(_07960_),
    .B2(\digitop_pav2.access_inst.access_ctrl0.state[14] ),
    .X(_10436_));
 a31o_1 _15229_ (.A1(net1319),
    .A2(_09524_),
    .A3(_09525_),
    .B1(_10436_),
    .X(_10437_));
 a31o_1 _15230_ (.A1(\digitop_pav2.access_inst.access_ctrl0.ld_dt_stb ),
    .A2(net1190),
    .A3(_10435_),
    .B1(_10437_),
    .X(_00019_));
 a21o_1 _15231_ (.A1(\digitop_pav2.access_inst.access_ctrl0.state[13] ),
    .A2(_09536_),
    .B1(_07397_),
    .X(_00018_));
 o21a_1 _15232_ (.A1(_07034_),
    .A2(net1210),
    .B1(\digitop_pav2.access_inst.access_check0.mem_sign_check_i ),
    .X(_10438_));
 o2111a_1 _15233_ (.A1(net1700),
    .A2(_07987_),
    .B1(_07970_),
    .C1(\digitop_pav2.access_inst.access_check0.mem_sign_check_sync_o ),
    .D1(net1235),
    .X(_10439_));
 a21o_1 _15234_ (.A1(\digitop_pav2.access_inst.access_ctrl0.rx_par1_i ),
    .A2(\digitop_pav2.access_inst.access_ctrl0.state[17] ),
    .B1(\digitop_pav2.access_inst.access_ctrl0.state[20] ),
    .X(_10440_));
 a31o_1 _15235_ (.A1(net1194),
    .A2(net818),
    .A3(_10440_),
    .B1(_10439_),
    .X(_10441_));
 or2_1 _15236_ (.A(_10438_),
    .B(_10441_),
    .X(_00017_));
 a32o_1 _15237_ (.A1(_07418_),
    .A2(_07480_),
    .A3(_10416_),
    .B1(net1206),
    .B2(net1145),
    .X(_10442_));
 a31o_1 _15238_ (.A1(\digitop_pav2.access_inst.access_check0.wr_lock_ck_i ),
    .A2(net1193),
    .A3(_08470_),
    .B1(_10442_),
    .X(_10443_));
 o21bai_1 _15239_ (.A1(_07505_),
    .A2(_10424_),
    .B1_N(_10443_),
    .Y(_00036_));
 a21o_1 _15240_ (.A1(\digitop_pav2.access_inst.access_ctrl0.ld_key_env_finish_i ),
    .A2(net366),
    .B1(net1201),
    .X(_10444_));
 a32o_1 _15241_ (.A1(\digitop_pav2.access_inst.access_ctrl0.ld_dt_stb ),
    .A2(net1190),
    .A3(_10434_),
    .B1(_10444_),
    .B2(net1144),
    .X(_00037_));
 or3b_1 _15242_ (.A(net1207),
    .B(net1235),
    .C_N(\digitop_pav2.access_inst.access_check0.pc_lock_check_sync_o ),
    .X(_10445_));
 a32o_1 _15243_ (.A1(net1258),
    .A2(net1319),
    .A3(_10416_),
    .B1(_10445_),
    .B2(\digitop_pav2.access_inst.access_check0.pc_lock_check_i ),
    .X(_10446_));
 a31o_1 _15244_ (.A1(\digitop_pav2.access_inst.access_check0.mem_sign_check_i ),
    .A2(_07321_),
    .A3(_09526_),
    .B1(_10446_),
    .X(_00038_));
 and3_1 _15245_ (.A(\digitop_pav2.ack_inst.state_ff[1] ),
    .B(net1248),
    .C(_08510_),
    .X(_10447_));
 a22o_1 _15246_ (.A1(\digitop_pav2.ack_inst.nvm_ack_rd_stb_o ),
    .A2(net1234),
    .B1(_10447_),
    .B2(_07062_),
    .X(_10448_));
 a31o_1 _15247_ (.A1(\digitop_pav2.ack_inst.state_ff[2] ),
    .A2(net1248),
    .A3(_07334_),
    .B1(_10448_),
    .X(_00042_));
 a32o_1 _15248_ (.A1(_09518_),
    .A2(_09521_),
    .A3(_10430_),
    .B1(_07960_),
    .B2(\digitop_pav2.access_inst.access_ctrl0.state[9] ),
    .X(_00039_));
 nor2_1 _15249_ (.A(net1188),
    .B(_09025_),
    .Y(_10449_));
 and3_1 _15250_ (.A(_07257_),
    .B(_07273_),
    .C(_09126_),
    .X(_10450_));
 a31o_1 _15251_ (.A1(net1293),
    .A2(net1197),
    .A3(_10450_),
    .B1(_10449_),
    .X(_00095_));
 or4_1 _15252_ (.A(net1186),
    .B(_07270_),
    .C(_07360_),
    .D(_09029_),
    .X(_10451_));
 and3_1 _15253_ (.A(net1294),
    .B(net1184),
    .C(_10451_),
    .X(_10452_));
 nor2_1 _15254_ (.A(_07364_),
    .B(_10451_),
    .Y(_10453_));
 a31o_1 _15255_ (.A1(net1295),
    .A2(net1195),
    .A3(_10453_),
    .B1(_10452_),
    .X(_00083_));
 nand2_2 _15256_ (.A(net1269),
    .B(_10398_),
    .Y(_10454_));
 inv_2 _15257_ (.A(_10454_),
    .Y(_10455_));
 nand2_1 _15258_ (.A(net1304),
    .B(_10454_),
    .Y(_10456_));
 o31a_1 _15259_ (.A1(net1296),
    .A2(net1249),
    .A3(_07273_),
    .B1(net1292),
    .X(_10457_));
 or2_2 _15260_ (.A(_07292_),
    .B(_09032_),
    .X(_10458_));
 inv_2 _15261_ (.A(_10458_),
    .Y(_10459_));
 or3_1 _15262_ (.A(net1195),
    .B(_07360_),
    .C(_10458_),
    .X(_10460_));
 nor3_1 _15263_ (.A(net1181),
    .B(_07271_),
    .C(_10460_),
    .Y(_10461_));
 nor2_1 _15264_ (.A(_07070_),
    .B(net1162),
    .Y(_10462_));
 nor2_1 _15265_ (.A(_09146_),
    .B(_09151_),
    .Y(_10463_));
 nand2_1 _15266_ (.A(net971),
    .B(\digitop_pav2.proc_ctrl_inst.ebv.state[2] ),
    .Y(_10464_));
 a21bo_1 _15267_ (.A1(net1303),
    .A2(_10464_),
    .B1_N(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[4] ),
    .X(_10465_));
 o21ba_1 _15268_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[12] ),
    .A2(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[3] ),
    .B1_N(net156),
    .X(_10466_));
 nor2_1 _15269_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.cg_en_13 ),
    .B(_10466_),
    .Y(_10467_));
 nand2_1 _15270_ (.A(_10465_),
    .B(_10467_),
    .Y(_10468_));
 o21a_1 _15271_ (.A1(net1296),
    .A2(net1251),
    .B1(net1291),
    .X(_10469_));
 o21a_1 _15272_ (.A1(net1188),
    .A2(_10456_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[11] ),
    .X(_10470_));
 o22a_1 _15273_ (.A1(net1290),
    .A2(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[9] ),
    .B1(net1188),
    .B2(net1296),
    .X(_10471_));
 nand2_1 _15274_ (.A(_07150_),
    .B(_10463_),
    .Y(_10472_));
 a221o_1 _15275_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[1] ),
    .A2(\digitop_pav2.proc_ctrl_inst.cmdfsm.pass_t1_i ),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdfsm.fm0x_dt_tx_st_i ),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[8] ),
    .C1(_10469_),
    .X(_10473_));
 a221o_1 _15276_ (.A1(net1290),
    .A2(net1195),
    .B1(_10472_),
    .B2(net1286),
    .C1(_10473_),
    .X(_10474_));
 or4_1 _15277_ (.A(_10462_),
    .B(_10468_),
    .C(_10471_),
    .D(_10474_),
    .X(_10475_));
 or4_4 _15278_ (.A(_08517_),
    .B(_10457_),
    .C(_10470_),
    .D(_10475_),
    .X(_10476_));
 inv_2 _15279_ (.A(_10476_),
    .Y(_10477_));
 nor2_1 _15280_ (.A(_07260_),
    .B(_09032_),
    .Y(_10478_));
 or3b_1 _15281_ (.A(_07291_),
    .B(_07331_),
    .C_N(_10478_),
    .X(_10479_));
 nor2_1 _15282_ (.A(net1181),
    .B(_10479_),
    .Y(_10480_));
 and3_1 _15283_ (.A(_07293_),
    .B(_07347_),
    .C(_10480_),
    .X(_10481_));
 a311o_1 _15284_ (.A1(net971),
    .A2(\digitop_pav2.proc_ctrl_inst.ebv.state[2] ),
    .A3(_07348_),
    .B1(_09027_),
    .C1(_10481_),
    .X(_10482_));
 a21oi_1 _15285_ (.A1(_07293_),
    .A2(_10476_),
    .B1(_10456_),
    .Y(_10483_));
 a22o_1 _15286_ (.A1(_10476_),
    .A2(_10482_),
    .B1(_10483_),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[11] ),
    .X(_00084_));
 a22o_1 _15287_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[12] ),
    .A2(net156),
    .B1(_08516_),
    .B2(_08518_),
    .X(_00085_));
 nand2_1 _15288_ (.A(net1217),
    .B(_08871_),
    .Y(_10484_));
 nor2_1 _15289_ (.A(_07087_),
    .B(_10484_),
    .Y(_10485_));
 a311o_1 _15290_ (.A1(net1287),
    .A2(_07315_),
    .A3(_09146_),
    .B1(_10485_),
    .C1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[1] ),
    .X(_10486_));
 and4_1 _15291_ (.A(net1287),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.pass_t1_i ),
    .C(_07301_),
    .D(_09146_),
    .X(_10487_));
 a31o_1 _15292_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.pass_t1_i ),
    .A2(_10476_),
    .A3(_10486_),
    .B1(_09142_),
    .X(_10488_));
 or2_1 _15293_ (.A(_10487_),
    .B(_10488_),
    .X(_00094_));
 a31o_1 _15294_ (.A1(_07330_),
    .A2(net1229),
    .A3(_10478_),
    .B1(_09018_),
    .X(_10489_));
 and2_1 _15295_ (.A(net1188),
    .B(_09024_),
    .X(_10490_));
 mux2_1 _15296_ (.A0(_09013_),
    .A1(_09024_),
    .S(net1188),
    .X(_10491_));
 nor2_1 _15297_ (.A(net1189),
    .B(_09020_),
    .Y(_10492_));
 a31o_1 _15298_ (.A1(_07290_),
    .A2(_07294_),
    .A3(_10489_),
    .B1(_10492_),
    .X(_10493_));
 o31a_1 _15299_ (.A1(_07367_),
    .A2(_10491_),
    .A3(_10493_),
    .B1(_10476_),
    .X(_10494_));
 and3_1 _15300_ (.A(net1293),
    .B(_07264_),
    .C(_10450_),
    .X(_10495_));
 a211o_1 _15301_ (.A1(net1290),
    .A2(_10477_),
    .B1(_10494_),
    .C1(_10495_),
    .X(_00093_));
 and2_1 _15302_ (.A(_07292_),
    .B(_07347_),
    .X(_10496_));
 a221o_1 _15303_ (.A1(net1189),
    .A2(_09021_),
    .B1(_10455_),
    .B2(_10496_),
    .C1(_09009_),
    .X(_10497_));
 nor2_1 _15304_ (.A(_07296_),
    .B(_09033_),
    .Y(_10498_));
 and3_1 _15305_ (.A(net1216),
    .B(_07283_),
    .C(_10498_),
    .X(_10499_));
 o2111a_1 _15306_ (.A1(net1184),
    .A2(_09126_),
    .B1(net1292),
    .C1(net1181),
    .D1(_07273_),
    .X(_10500_));
 a22o_1 _15307_ (.A1(_07048_),
    .A2(_07298_),
    .B1(_10476_),
    .B2(_10497_),
    .X(_10501_));
 a211o_1 _15308_ (.A1(net1291),
    .A2(_10477_),
    .B1(_10499_),
    .C1(_10501_),
    .X(_10502_));
 a31o_1 _15309_ (.A1(net1293),
    .A2(net1198),
    .A3(_09127_),
    .B1(_10500_),
    .X(_10503_));
 or2_1 _15310_ (.A(_10502_),
    .B(_10503_),
    .X(_00092_));
 or2_1 _15311_ (.A(net1162),
    .B(_10477_),
    .X(_10504_));
 and2_2 _15312_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[5] ),
    .B(_07331_),
    .X(_10505_));
 nor2_1 _15313_ (.A(_08518_),
    .B(_10505_),
    .Y(_10506_));
 a2bb2o_1 _15314_ (.A1_N(_08516_),
    .A2_N(_10506_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[8] ),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.fm0x_dt_tx_st_i ),
    .X(_10507_));
 a22o_1 _15315_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[5] ),
    .A2(_10504_),
    .B1(_10507_),
    .B2(_10476_),
    .X(_00091_));
 and2_1 _15316_ (.A(_07348_),
    .B(_10464_),
    .X(_10508_));
 a31o_1 _15317_ (.A1(_07295_),
    .A2(net1229),
    .A3(net1188),
    .B1(_10508_),
    .X(_00090_));
 a22o_1 _15318_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[3] ),
    .A2(net156),
    .B1(_08516_),
    .B2(_10505_),
    .X(_00089_));
 a21o_1 _15319_ (.A1(net1181),
    .A2(_07274_),
    .B1(_10504_),
    .X(_10509_));
 nor2_1 _15320_ (.A(_07244_),
    .B(_07279_),
    .Y(_10510_));
 and2b_1 _15321_ (.A_N(net1249),
    .B(_10510_),
    .X(_10511_));
 and2b_1 _15322_ (.A_N(_09127_),
    .B(_10511_),
    .X(_10512_));
 and2_1 _15323_ (.A(_07270_),
    .B(_07365_),
    .X(_10513_));
 and3_1 _15324_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[11] ),
    .B(net1181),
    .C(net1188),
    .X(_10514_));
 a211o_1 _15325_ (.A1(net1304),
    .A2(_10514_),
    .B1(_10513_),
    .C1(_07326_),
    .X(_10515_));
 o31a_1 _15326_ (.A1(net1198),
    .A2(_07264_),
    .A3(net1197),
    .B1(net1292),
    .X(_10516_));
 a311o_1 _15327_ (.A1(_07274_),
    .A2(_07276_),
    .A3(_10516_),
    .B1(_10515_),
    .C1(_10512_),
    .X(_10517_));
 a22o_1 _15328_ (.A1(_07278_),
    .A2(_10509_),
    .B1(_10517_),
    .B2(_10476_),
    .X(_00088_));
 o22a_1 _15329_ (.A1(_07150_),
    .A2(_10477_),
    .B1(_10485_),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[1] ),
    .X(_10518_));
 a41o_1 _15330_ (.A1(net1287),
    .A2(_07150_),
    .A3(_07316_),
    .A4(_09146_),
    .B1(_10518_),
    .X(_00087_));
 nor2_1 _15331_ (.A(_07274_),
    .B(_09126_),
    .Y(_10519_));
 a31o_1 _15332_ (.A1(net1292),
    .A2(net1181),
    .A3(_07325_),
    .B1(_10516_),
    .X(_10520_));
 o21a_1 _15333_ (.A1(_07277_),
    .A2(_10460_),
    .B1(net1292),
    .X(_10521_));
 and2_1 _15334_ (.A(net1289),
    .B(net1197),
    .X(_10522_));
 or2_2 _15335_ (.A(_07318_),
    .B(_10522_),
    .X(_10523_));
 and3b_1 _15336_ (.A_N(_09158_),
    .B(_07298_),
    .C(net1251),
    .X(_10524_));
 and3_1 _15337_ (.A(net1294),
    .B(_07311_),
    .C(_10453_),
    .X(_10525_));
 a221o_1 _15338_ (.A1(_09152_),
    .A2(_10523_),
    .B1(_10525_),
    .B2(_07248_),
    .C1(_10524_),
    .X(_10526_));
 and4_1 _15339_ (.A(net1251),
    .B(_07296_),
    .C(net1183),
    .D(_09158_),
    .X(_10527_));
 o21a_1 _15340_ (.A1(_09033_),
    .A2(_10527_),
    .B1(_07283_),
    .X(_10528_));
 a2bb2o_1 _15341_ (.A1_N(_10478_),
    .A2_N(_07352_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[5] ),
    .B2(_10458_),
    .X(_10529_));
 nand2_1 _15342_ (.A(net1249),
    .B(net1186),
    .Y(_10530_));
 and3_1 _15343_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.piex_dt_rx_done ),
    .B(net1293),
    .C(net1186),
    .X(_10531_));
 and3_1 _15344_ (.A(net1251),
    .B(_07284_),
    .C(_09130_),
    .X(_10532_));
 or2_1 _15345_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[9] ),
    .B(_07350_),
    .X(_10533_));
 o21a_1 _15346_ (.A1(net1290),
    .A2(_10533_),
    .B1(net1296),
    .X(_10534_));
 or3b_1 _15347_ (.A(_10534_),
    .B(_09176_),
    .C_N(_10467_),
    .X(_10535_));
 a32o_1 _15348_ (.A1(_07328_),
    .A2(_08870_),
    .A3(_09151_),
    .B1(_09032_),
    .B2(net1286),
    .X(_10536_));
 or4_1 _15349_ (.A(_10531_),
    .B(_10532_),
    .C(_10535_),
    .D(_10536_),
    .X(_10537_));
 and3_1 _15350_ (.A(_07293_),
    .B(_07347_),
    .C(_10479_),
    .X(_10538_));
 and3_1 _15351_ (.A(_07290_),
    .B(_07330_),
    .C(_07363_),
    .X(_10539_));
 a31o_1 _15352_ (.A1(_07261_),
    .A2(_07293_),
    .A3(_10539_),
    .B1(_10538_),
    .X(_10540_));
 or4_1 _15353_ (.A(_10528_),
    .B(_10529_),
    .C(_10537_),
    .D(_10540_),
    .X(_10541_));
 a2111o_1 _15354_ (.A1(_10519_),
    .A2(_10520_),
    .B1(_10521_),
    .C1(_10526_),
    .D1(_10541_),
    .X(_10542_));
 mux2_1 _15355_ (.A0(net1294),
    .A1(_10542_),
    .S(_10476_),
    .X(_00082_));
 a22o_1 _15356_ (.A1(_07111_),
    .A2(\digitop_pav2.proc_ctrl_inst.ebv.state[4] ),
    .B1(_09664_),
    .B2(_07071_),
    .X(_00096_));
 or3_1 _15357_ (.A(_07329_),
    .B(_08871_),
    .C(_09151_),
    .X(_10543_));
 a31o_1 _15358_ (.A1(net1304),
    .A2(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[7] ),
    .A3(net1195),
    .B1(_09141_),
    .X(_10544_));
 nand2_1 _15359_ (.A(net1288),
    .B(_07300_),
    .Y(_10545_));
 o21ai_1 _15360_ (.A1(_07300_),
    .A2(_07302_),
    .B1(net1287),
    .Y(_10546_));
 nor2_1 _15361_ (.A(_09146_),
    .B(_10546_),
    .Y(_10547_));
 or3b_1 _15362_ (.A(_10544_),
    .B(_10547_),
    .C_N(_10543_),
    .X(_10548_));
 a221o_1 _15363_ (.A1(net1286),
    .A2(_10461_),
    .B1(_10463_),
    .B2(_10523_),
    .C1(_10548_),
    .X(_10549_));
 or3_1 _15364_ (.A(_09128_),
    .B(_09140_),
    .C(_10549_),
    .X(_10550_));
 mux2_1 _15365_ (.A0(net1286),
    .A1(_10550_),
    .S(_10476_),
    .X(_00086_));
 a31o_1 _15366_ (.A1(_07032_),
    .A2(_07033_),
    .A3(_07417_),
    .B1(_07576_),
    .X(_10551_));
 mux2_1 _15367_ (.A0(\digitop_pav2.access_inst.access_ctrl0.state[23] ),
    .A1(\digitop_pav2.access_inst.access_ctrl0.state[10] ),
    .S(_07960_),
    .X(_10552_));
 a41o_1 _15368_ (.A1(\digitop_pav2.access_inst.access_check0.pc_lock_check_sync_o ),
    .A2(\digitop_pav2.access_inst.access_check0.pc_lock_check_i ),
    .A3(_09521_),
    .A4(_10426_),
    .B1(_10552_),
    .X(_10553_));
 a31o_1 _15369_ (.A1(_08470_),
    .A2(_09525_),
    .A3(_10551_),
    .B1(_10553_),
    .X(_10554_));
 a31o_1 _15370_ (.A1(_07024_),
    .A2(net1145),
    .A3(net1191),
    .B1(_10554_),
    .X(_00015_));
 and2_1 _15371_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[6] ),
    .B(_10326_),
    .X(_10555_));
 or4_1 _15372_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[6] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[5] ),
    .C(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[0] ),
    .D(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[7] ),
    .X(_10556_));
 or4_1 _15373_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[4] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[3] ),
    .C(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[2] ),
    .D(_10556_),
    .X(_10557_));
 o21a_1 _15374_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[1] ),
    .A2(_10557_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.state[2] ),
    .X(_10558_));
 and4b_1 _15375_ (.A_N(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[6] ),
    .B(_10410_),
    .C(_10411_),
    .D(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[5] ),
    .X(_10559_));
 a22o_1 _15376_ (.A1(_07909_),
    .A2(_10413_),
    .B1(_10559_),
    .B2(_07900_),
    .X(_10560_));
 and2_1 _15377_ (.A(_10344_),
    .B(_10560_),
    .X(_10561_));
 a31o_1 _15378_ (.A1(_10399_),
    .A2(_10558_),
    .A3(_10561_),
    .B1(_10555_),
    .X(_00074_));
 and3_1 _15379_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[7] ),
    .B(_07861_),
    .C(_07867_),
    .X(_10562_));
 a32o_1 _15380_ (.A1(_10399_),
    .A2(_10413_),
    .A3(_10562_),
    .B1(_10326_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.state[5] ),
    .X(_00073_));
 or4b_1 _15381_ (.A(_10333_),
    .B(_10337_),
    .C(_10335_),
    .D_N(\digitop_pav2.invent_inst.invent_sel_pav2.state[0] ),
    .X(_10563_));
 a2bb2o_1 _15382_ (.A1_N(_10346_),
    .A2_N(_10563_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.state[4] ),
    .B2(_10326_),
    .X(_00072_));
 or3_1 _15383_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[6] ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.state[7] ),
    .C(_10328_),
    .X(_10564_));
 or2_1 _15384_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[2] ),
    .B(_10564_),
    .X(_10565_));
 inv_2 _15385_ (.A(_10565_),
    .Y(_10566_));
 nand2b_1 _15386_ (.A_N(net1173),
    .B(net1174),
    .Y(_10567_));
 or2_1 _15387_ (.A(net1175),
    .B(_10567_),
    .X(_10568_));
 nor2_1 _15388_ (.A(_10400_),
    .B(_10567_),
    .Y(_10569_));
 nand2_2 _15389_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[0] ),
    .B(net1175),
    .Y(_10570_));
 and4_2 _15390_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[0] ),
    .B(net1175),
    .C(net1174),
    .D(net1173),
    .X(_10571_));
 nor2_1 _15391_ (.A(_10567_),
    .B(_10570_),
    .Y(_10572_));
 nor2_1 _15392_ (.A(_10401_),
    .B(_10408_),
    .Y(_10573_));
 or2_1 _15393_ (.A(_10401_),
    .B(_10408_),
    .X(_10574_));
 and4b_1 _15394_ (.A_N(net1175),
    .B(net1174),
    .C(net1173),
    .D(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[0] ),
    .X(_10575_));
 a221o_1 _15395_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[9] ),
    .A2(_10572_),
    .B1(_10575_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[3] ),
    .C1(_10573_),
    .X(_10576_));
 a221o_1 _15396_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[12] ),
    .A2(_10569_),
    .B1(_10571_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[1] ),
    .C1(_10576_),
    .X(_10577_));
 nand2_1 _15397_ (.A(_07137_),
    .B(net1175),
    .Y(_10578_));
 and4_1 _15398_ (.A(_07137_),
    .B(net1175),
    .C(net1174),
    .D(net1173),
    .X(_10579_));
 and4bb_1 _15399_ (.A_N(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[0] ),
    .B_N(net1175),
    .C(net1174),
    .D(net1173),
    .X(_10580_));
 a22o_1 _15400_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[2] ),
    .A2(_10579_),
    .B1(_10580_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[4] ),
    .X(_10581_));
 nor2_1 _15401_ (.A(_10567_),
    .B(_10578_),
    .Y(_10582_));
 nor2_1 _15402_ (.A(_10409_),
    .B(_10578_),
    .Y(_10583_));
 a22o_1 _15403_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[10] ),
    .A2(_10582_),
    .B1(_10583_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[6] ),
    .X(_10584_));
 nor2_1 _15404_ (.A(_10408_),
    .B(_10567_),
    .Y(_10585_));
 a221o_1 _15405_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[0] ),
    .A2(_10402_),
    .B1(_10585_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[11] ),
    .C1(_10584_),
    .X(_10586_));
 nor2_1 _15406_ (.A(_10401_),
    .B(_10578_),
    .Y(_10587_));
 nor2_1 _15407_ (.A(_10401_),
    .B(_10570_),
    .Y(_10588_));
 nor2_2 _15408_ (.A(_10409_),
    .B(_10570_),
    .Y(_10589_));
 nor2_1 _15409_ (.A(_10400_),
    .B(_10409_),
    .Y(_10590_));
 a22o_1 _15410_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[5] ),
    .A2(_10589_),
    .B1(_10590_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[8] ),
    .X(_10591_));
 a221o_1 _15411_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[14] ),
    .A2(_10587_),
    .B1(_10588_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[13] ),
    .C1(_10591_),
    .X(_10592_));
 a2111o_1 _15412_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[7] ),
    .A2(_10410_),
    .B1(_10581_),
    .C1(_10586_),
    .D1(_10592_),
    .X(_10593_));
 nor2_1 _15413_ (.A(_10577_),
    .B(_10593_),
    .Y(_10594_));
 xor2_1 _15414_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[5] ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[6] ),
    .X(_10595_));
 nand2_1 _15415_ (.A(_10411_),
    .B(_10595_),
    .Y(_10596_));
 nor2_1 _15416_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[15] ),
    .B(_10574_),
    .Y(_10597_));
 a221o_1 _15417_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[12] ),
    .A2(_10569_),
    .B1(_10585_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[11] ),
    .C1(_10573_),
    .X(_10598_));
 a221o_1 _15418_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[1] ),
    .A2(_10571_),
    .B1(_10572_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[9] ),
    .C1(_10598_),
    .X(_10599_));
 a22o_1 _15419_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[3] ),
    .A2(_10575_),
    .B1(_10588_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[13] ),
    .X(_10600_));
 a22o_1 _15420_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[4] ),
    .A2(_10580_),
    .B1(_10582_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[10] ),
    .X(_10601_));
 a221o_1 _15421_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[7] ),
    .A2(_10410_),
    .B1(_10579_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[2] ),
    .C1(_10601_),
    .X(_10602_));
 a22o_1 _15422_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[0] ),
    .A2(_10402_),
    .B1(_10589_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[5] ),
    .X(_10603_));
 a221o_1 _15423_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[14] ),
    .A2(_10587_),
    .B1(_10590_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[8] ),
    .C1(_10603_),
    .X(_10604_));
 a2111o_1 _15424_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[6] ),
    .A2(_10583_),
    .B1(_10600_),
    .C1(_10602_),
    .D1(_10604_),
    .X(_10605_));
 nor2_1 _15425_ (.A(_10599_),
    .B(_10605_),
    .Y(_10606_));
 o21ai_1 _15426_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[15] ),
    .A2(_10574_),
    .B1(_10596_),
    .Y(_10607_));
 o32a_1 _15427_ (.A1(_10594_),
    .A2(_10596_),
    .A3(_10597_),
    .B1(_10606_),
    .B2(_10607_),
    .X(_10608_));
 xor2_1 _15428_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[7] ),
    .B(_10608_),
    .X(_10609_));
 mux2_1 _15429_ (.A0(_10405_),
    .A1(_10411_),
    .S(_10407_),
    .X(_10610_));
 nand2_1 _15430_ (.A(_10609_),
    .B(_10610_),
    .Y(_10611_));
 xnor2_1 _15431_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[7] ),
    .B(_10568_),
    .Y(_10612_));
 or4bb_1 _15432_ (.A(_10411_),
    .B(_10612_),
    .C_N(_10405_),
    .D_N(_10407_),
    .X(_10613_));
 nor2_1 _15433_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[4] ),
    .B(_10574_),
    .Y(_10614_));
 a221o_1 _15434_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[4] ),
    .A2(_10580_),
    .B1(_10588_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[13] ),
    .C1(_10411_),
    .X(_10615_));
 a221o_1 _15435_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[12] ),
    .A2(_10569_),
    .B1(_10572_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[9] ),
    .C1(_10615_),
    .X(_10616_));
 a22o_1 _15436_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[0] ),
    .A2(_10402_),
    .B1(_10575_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[3] ),
    .X(_10617_));
 a22o_1 _15437_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[6] ),
    .A2(_10583_),
    .B1(_10590_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[8] ),
    .X(_10618_));
 a221o_1 _15438_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[10] ),
    .A2(_10582_),
    .B1(_10585_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[11] ),
    .C1(_10618_),
    .X(_10619_));
 a22o_1 _15439_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[2] ),
    .A2(_10579_),
    .B1(_10589_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[5] ),
    .X(_10620_));
 a221o_1 _15440_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[7] ),
    .A2(_10410_),
    .B1(_10573_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[15] ),
    .C1(_10620_),
    .X(_10621_));
 a2111o_1 _15441_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[14] ),
    .A2(_10587_),
    .B1(_10617_),
    .C1(_10619_),
    .D1(_10621_),
    .X(_10622_));
 and2_1 _15442_ (.A(\digitop_pav2.boot_inst.boot_proc0.proc_mask[17] ),
    .B(_10571_),
    .X(_10623_));
 a22o_1 _15443_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[22] ),
    .A2(_10583_),
    .B1(_10589_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[21] ),
    .X(_10624_));
 a221o_1 _15444_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[20] ),
    .A2(_10580_),
    .B1(_10588_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[29] ),
    .C1(_10624_),
    .X(_10625_));
 a22o_1 _15445_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[25] ),
    .A2(_10572_),
    .B1(_10582_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[26] ),
    .X(_10626_));
 a22o_1 _15446_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[28] ),
    .A2(_10569_),
    .B1(_10585_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[27] ),
    .X(_10627_));
 or4b_1 _15447_ (.A(_10623_),
    .B(_10626_),
    .C(_10627_),
    .D_N(_10411_),
    .X(_10628_));
 a221o_1 _15448_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[16] ),
    .A2(_10402_),
    .B1(_10590_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[24] ),
    .C1(_10628_),
    .X(_10629_));
 a22o_1 _15449_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[19] ),
    .A2(_10575_),
    .B1(_10579_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[18] ),
    .X(_10630_));
 a221o_1 _15450_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[23] ),
    .A2(_10410_),
    .B1(_10587_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[30] ),
    .C1(_10630_),
    .X(_10631_));
 or3_1 _15451_ (.A(_10625_),
    .B(_10629_),
    .C(_10631_),
    .X(_10632_));
 o21a_1 _15452_ (.A1(_10616_),
    .A2(_10622_),
    .B1(_10632_),
    .X(_10633_));
 and2_1 _15453_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[4] ),
    .B(_10571_),
    .X(_10634_));
 a221o_1 _15454_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[31] ),
    .A2(_10614_),
    .B1(_10634_),
    .B2(\digitop_pav2.boot_inst.boot_proc0.proc_mask[1] ),
    .C1(_10633_),
    .X(_10635_));
 xor2_1 _15455_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[7] ),
    .B(_10635_),
    .X(_10636_));
 a32o_1 _15456_ (.A1(_10344_),
    .A2(_10611_),
    .A3(_10613_),
    .B1(_10636_),
    .B2(_10337_),
    .X(_10637_));
 a21o_1 _15457_ (.A1(_10565_),
    .A2(_10637_),
    .B1(_10345_),
    .X(_10638_));
 and4_1 _15458_ (.A(_10382_),
    .B(_10383_),
    .C(_10386_),
    .D(_10388_),
    .X(_10639_));
 or4bb_1 _15459_ (.A(_10373_),
    .B(_10375_),
    .C_N(_10380_),
    .D_N(_10639_),
    .X(_10640_));
 o31a_1 _15460_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[1] ),
    .A2(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[0] ),
    .A3(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[7] ),
    .B1(_10557_),
    .X(_10641_));
 a2111o_1 _15461_ (.A1(_10378_),
    .A2(_10640_),
    .B1(_10641_),
    .C1(_07860_),
    .D1(_07858_),
    .X(_10642_));
 nor2_1 _15462_ (.A(_10376_),
    .B(_10380_),
    .Y(_10643_));
 mux2_1 _15463_ (.A0(_10372_),
    .A1(_10639_),
    .S(_10643_),
    .X(_10644_));
 a21bo_1 _15464_ (.A1(_10375_),
    .A2(_10378_),
    .B1_N(_07869_),
    .X(_10645_));
 or3b_1 _15465_ (.A(_10645_),
    .B(_10373_),
    .C_N(_10644_),
    .X(_10646_));
 a22o_1 _15466_ (.A1(_10337_),
    .A2(_10642_),
    .B1(_10646_),
    .B2(_10344_),
    .X(_10647_));
 a31o_1 _15467_ (.A1(_10341_),
    .A2(_10566_),
    .A3(_10647_),
    .B1(_10638_),
    .X(_10648_));
 inv_2 _15468_ (.A(_10648_),
    .Y(_10649_));
 and4_1 _15469_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[9] ),
    .B(_10325_),
    .C(_10341_),
    .D(_10648_),
    .X(_10650_));
 or3b_1 _15470_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[1] ),
    .B(_10557_),
    .C_N(\digitop_pav2.invent_inst.invent_sel_pav2.state[2] ),
    .X(_10651_));
 nand2_1 _15471_ (.A(_07128_),
    .B(_10651_),
    .Y(_10652_));
 a32o_1 _15472_ (.A1(net1014),
    .A2(_10565_),
    .A3(_10652_),
    .B1(_10331_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.select_valid_o ),
    .X(_10653_));
 o211a_1 _15473_ (.A1(_10558_),
    .A2(_10564_),
    .B1(_07128_),
    .C1(_10325_),
    .X(_10654_));
 a211o_1 _15474_ (.A1(_10398_),
    .A2(_10654_),
    .B1(_10653_),
    .C1(_10650_),
    .X(_00071_));
 and4_1 _15475_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[9] ),
    .B(net1014),
    .C(_10341_),
    .D(_10649_),
    .X(_10655_));
 and3b_1 _15476_ (.A_N(_10561_),
    .B(_10558_),
    .C(_10399_),
    .X(_10656_));
 a211o_1 _15477_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[2] ),
    .A2(_10326_),
    .B1(_10655_),
    .C1(_10656_),
    .X(_00070_));
 a22o_1 _15478_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[1] ),
    .A2(_10326_),
    .B1(_10328_),
    .B2(_10399_),
    .X(_00069_));
 o31a_1 _15479_ (.A1(_10326_),
    .A2(_10333_),
    .A3(_10335_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.state[0] ),
    .X(_00064_));
 mux2_1 _15480_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_i ),
    .A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_s_ff_i ),
    .S(\digitop_pav2.invent_inst.invent_qqqr_pav2.query_inversion ),
    .X(_10657_));
 xnor2_1 _15481_ (.A(net1178),
    .B(_10657_),
    .Y(_10658_));
 xnor2_1 _15482_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.s1_i ),
    .B(net1178),
    .Y(_10659_));
 xnor2_1 _15483_ (.A(net1178),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ),
    .Y(_10660_));
 xnor2_1 _15484_ (.A(net1178),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.s0_i ),
    .Y(_10661_));
 o21ai_1 _15485_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[5] ),
    .A2(\digitop_pav2.invent_inst.invent_qqqr_pav2.sl_i ),
    .B1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[4] ),
    .Y(_10662_));
 a21o_1 _15486_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[5] ),
    .A2(\digitop_pav2.invent_inst.invent_qqqr_pav2.sl_i ),
    .B1(_10662_),
    .X(_10663_));
 xnor2_1 _15487_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_s_ff_i ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[0] ),
    .Y(_10664_));
 and4b_1 _15488_ (.A_N(\digitop_pav2.invent_inst.invent_qqqr_pav2.query_inversion ),
    .B(_10660_),
    .C(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[7] ),
    .D(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[6] ),
    .X(_10665_));
 a31o_1 _15489_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[7] ),
    .A2(_07133_),
    .A3(_10659_),
    .B1(_10665_),
    .X(_10666_));
 and4_1 _15490_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[7] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[6] ),
    .C(\digitop_pav2.invent_inst.invent_qqqr_pav2.query_inversion ),
    .D(_10664_),
    .X(_10667_));
 a311o_1 _15491_ (.A1(_07132_),
    .A2(_07133_),
    .A3(_10661_),
    .B1(_10666_),
    .C1(_10667_),
    .X(_10668_));
 a31o_1 _15492_ (.A1(_07132_),
    .A2(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[6] ),
    .A3(_10658_),
    .B1(_10668_),
    .X(_10669_));
 nand2_1 _15493_ (.A(_10663_),
    .B(_10669_),
    .Y(_10670_));
 xor2_1 _15494_ (.A(\digitop_pav2.dr ),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[1] ),
    .X(_10671_));
 nand2_1 _15495_ (.A(net1180),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[0] ),
    .Y(_10672_));
 or2_1 _15496_ (.A(net1180),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[0] ),
    .X(_10673_));
 a21oi_1 _15497_ (.A1(_10672_),
    .A2(_10673_),
    .B1(_10671_),
    .Y(_10674_));
 xnor2_1 _15498_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[3] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[4] ),
    .Y(_10675_));
 nand2_1 _15499_ (.A(net1179),
    .B(_08975_),
    .Y(_10676_));
 o211ai_1 _15500_ (.A1(net1179),
    .A2(_10675_),
    .B1(_10676_),
    .C1(_10674_),
    .Y(_10677_));
 and3_1 _15501_ (.A(net1277),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[0] ),
    .C(_07238_),
    .X(_10678_));
 and4bb_1 _15502_ (.A_N(net1282),
    .B_N(_10674_),
    .C(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[0] ),
    .D(net1279),
    .X(_10679_));
 a221o_1 _15503_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[7] ),
    .A2(_10670_),
    .B1(_10677_),
    .B2(_10678_),
    .C1(_10679_),
    .X(_10680_));
 a21o_1 _15504_ (.A1(_07336_),
    .A2(_10680_),
    .B1(\digitop_pav2.invent_inst.invent_qqqr_pav2.r_invent3_o ),
    .X(_00057_));
 a31o_1 _15505_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[7] ),
    .A2(_10663_),
    .A3(_10669_),
    .B1(net808),
    .X(_10681_));
 o22a_1 _15506_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[11] ),
    .A2(_07336_),
    .B1(_10681_),
    .B2(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[4] ),
    .X(_00056_));
 or2_1 _15507_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[0] ),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[1] ),
    .X(_10682_));
 or4_1 _15508_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[2] ),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[3] ),
    .C(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[4] ),
    .D(_10682_),
    .X(_10683_));
 or3_2 _15509_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[5] ),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[6] ),
    .C(_10683_),
    .X(_10684_));
 inv_2 _15510_ (.A(_10684_),
    .Y(_10685_));
 or3_1 _15511_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[7] ),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[8] ),
    .C(_10684_),
    .X(_10686_));
 or2_1 _15512_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[9] ),
    .B(_10686_),
    .X(_10687_));
 or3_1 _15513_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[10] ),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[11] ),
    .C(_10687_),
    .X(_10688_));
 or2_1 _15514_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[12] ),
    .B(_10688_),
    .X(_10689_));
 nor2_1 _15515_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[13] ),
    .B(_10689_),
    .Y(_10690_));
 and2b_1 _15516_ (.A_N(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[14] ),
    .B(_10690_),
    .X(_10691_));
 or2_1 _15517_ (.A(_07244_),
    .B(net1225),
    .X(_10692_));
 or2_1 _15518_ (.A(net1247),
    .B(_10692_),
    .X(_10693_));
 nor2_1 _15519_ (.A(\digitop_pav2.proc_ctrl_inst.int_timeout_t2 ),
    .B(_10693_),
    .Y(_10694_));
 and2b_2 _15520_ (.A_N(net1722),
    .B(net1713),
    .X(_10695_));
 nand2b_1 _15521_ (.A_N(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[2] ),
    .B(net1713),
    .Y(_10696_));
 or2_1 _15522_ (.A(net1718),
    .B(net1714),
    .X(_10697_));
 inv_2 _15523_ (.A(_10697_),
    .Y(_10698_));
 nand4b_1 _15524_ (.A_N(net1282),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[0] ),
    .C(_10674_),
    .D(net1279),
    .Y(_10699_));
 o32a_1 _15525_ (.A1(_10694_),
    .A2(net1719),
    .A3(_10699_),
    .B1(_07127_),
    .B2(net1677),
    .X(_10700_));
 o21ai_1 _15526_ (.A1(_07020_),
    .A2(_10691_),
    .B1(net1720),
    .Y(_10701_));
 a21o_1 _15527_ (.A1(_07336_),
    .A2(_10701_),
    .B1(\digitop_pav2.invent_inst.invent_qqqr_pav2.r_invent2_o ),
    .X(_00055_));
 a2bb2o_1 _15528_ (.A1_N(_10694_),
    .A2_N(_10697_),
    .B1(net1714),
    .B2(_09097_),
    .X(_10702_));
 nand2b_1 _15529_ (.A_N(_10677_),
    .B(_10678_),
    .Y(_10703_));
 or2_1 _15530_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[1] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[6] ),
    .X(_10704_));
 nand2_1 _15531_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[1] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[6] ),
    .Y(_10705_));
 nand2_1 _15532_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[0] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[7] ),
    .Y(_10706_));
 or2_1 _15533_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[0] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[7] ),
    .X(_10707_));
 a22o_1 _15534_ (.A1(_10704_),
    .A2(_10705_),
    .B1(_10706_),
    .B2(_10707_),
    .X(_10708_));
 and4b_1 _15535_ (.A_N(net1672),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[0] ),
    .C(_07238_),
    .D(net1274),
    .X(_10709_));
 nand2b_1 _15536_ (.A_N(_10708_),
    .B(_10709_),
    .Y(_10710_));
 a31o_1 _15537_ (.A1(_10699_),
    .A2(_10703_),
    .A3(_10710_),
    .B1(net808),
    .X(_10711_));
 a2bb2o_1 _15538_ (.A1_N(net1715),
    .A2_N(_10711_),
    .B1(\digitop_pav2.invent_inst.invent_qqqr_pav2.flags_en_o ),
    .B2(net808),
    .X(_00063_));
 or2_1 _15539_ (.A(net1715),
    .B(_10708_),
    .X(_10712_));
 a221o_1 _15540_ (.A1(net1677),
    .A2(\digitop_pav2.invent_inst.invent_qqqr_pav2.flags_en_o ),
    .B1(_10709_),
    .B2(net1716),
    .C1(net808),
    .X(_10713_));
 o21a_1 _15541_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[7] ),
    .A2(_07336_),
    .B1(_10713_),
    .X(_00062_));
 a221o_1 _15542_ (.A1(net1675),
    .A2(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[0] ),
    .B1(_10691_),
    .B2(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[3] ),
    .C1(net808),
    .X(_10714_));
 o21a_1 _15543_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[6] ),
    .A2(_07336_),
    .B1(_10714_),
    .X(_00061_));
 a32o_1 _15544_ (.A1(net1144),
    .A2(net1190),
    .A3(_07524_),
    .B1(_07960_),
    .B2(\digitop_pav2.access_inst.access_ctrl0.state[11] ),
    .X(_10715_));
 a31o_1 _15545_ (.A1(net1148),
    .A2(net1190),
    .A3(_08470_),
    .B1(_10715_),
    .X(_00016_));
 nor2_1 _15546_ (.A(net808),
    .B(_10703_),
    .Y(_10716_));
 a22o_1 _15547_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[4] ),
    .A2(net808),
    .B1(net1715),
    .B2(_10716_),
    .X(_00060_));
 or4_1 _15548_ (.A(_07337_),
    .B(_09096_),
    .C(_10695_),
    .D(_10699_),
    .X(_10717_));
 a21bo_1 _15549_ (.A1(net1172),
    .A2(_07337_),
    .B1_N(_10717_),
    .X(_00059_));
 a31o_1 _15550_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[5] ),
    .A2(_07336_),
    .A3(net1165),
    .B1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[1] ),
    .X(_00058_));
 and2_1 _15551_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[0] ),
    .B(net808),
    .X(_00054_));
 nand2_1 _15552_ (.A(net1445),
    .B(net159),
    .Y(_10718_));
 and2_1 _15553_ (.A(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_crc_en ),
    .B(net1431),
    .X(_10719_));
 nand2_1 _15554_ (.A(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_crc_en ),
    .B(net1431),
    .Y(_10720_));
 nor2_1 _15555_ (.A(_07058_),
    .B(_10720_),
    .Y(_10721_));
 a41o_1 _15556_ (.A1(\digitop_pav2.boot_inst.boot_ctrl0.state[2] ),
    .A2(net1432),
    .A3(net159),
    .A4(_07836_),
    .B1(_10721_),
    .X(_10722_));
 a21o_1 _15557_ (.A1(_07058_),
    .A2(_07837_),
    .B1(_07059_),
    .X(_10723_));
 nand2_1 _15558_ (.A(net1431),
    .B(_10723_),
    .Y(_10724_));
 a21o_1 _15559_ (.A1(\digitop_pav2.boot_inst.boot_ctrl0.state[3] ),
    .A2(_10724_),
    .B1(_10722_),
    .X(_00053_));
 a21oi_1 _15560_ (.A1(_07059_),
    .A2(\digitop_pav2.boot_inst.boot_ctrl0.state[3] ),
    .B1(\digitop_pav2.boot_inst.boot_ctrl0.state[0] ),
    .Y(_10725_));
 nand2_1 _15561_ (.A(_07058_),
    .B(net1321),
    .Y(_10726_));
 o2bb2a_1 _15562_ (.A1_N(\digitop_pav2.boot_inst.boot_ctrl0.state[2] ),
    .A2_N(_10718_),
    .B1(_10725_),
    .B2(net1400),
    .X(_10727_));
 nand2_1 _15563_ (.A(_10726_),
    .B(_10727_),
    .Y(_00052_));
 and3_1 _15564_ (.A(\digitop_pav2.boot_inst.boot_ctrl0.proc_boot_end_i ),
    .B(net1431),
    .C(\digitop_pav2.boot_inst.boot_ctrl0.state[3] ),
    .X(_10728_));
 nor2_1 _15565_ (.A(_07836_),
    .B(_10718_),
    .Y(_10729_));
 a32o_1 _15566_ (.A1(_07058_),
    .A2(_07837_),
    .A3(_10728_),
    .B1(net1400),
    .B2(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_crc_en ),
    .X(_10730_));
 a21o_1 _15567_ (.A1(\digitop_pav2.boot_inst.boot_ctrl0.state[2] ),
    .A2(_10729_),
    .B1(_10730_),
    .X(_00051_));
 xnor2_1 _15568_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[0] ),
    .B(_08896_),
    .Y(_10731_));
 xnor2_2 _15569_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[0] ),
    .B(_08895_),
    .Y(_10732_));
 and3_1 _15570_ (.A(net470),
    .B(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_2b_o ),
    .C(_10732_),
    .X(_10733_));
 and4b_1 _15571_ (.A_N(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[2] ),
    .B(_07040_),
    .C(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[0] ),
    .D(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[3] ),
    .X(_10734_));
 or4bb_1 _15572_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[1] ),
    .C_N(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[0] ),
    .D_N(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[3] ),
    .X(_10735_));
 o211a_1 _15573_ (.A1(_10731_),
    .A2(_10734_),
    .B1(net463),
    .C1(net413),
    .X(_10736_));
 a211o_1 _15574_ (.A1(net426),
    .A2(_07112_),
    .B1(_10733_),
    .C1(_10736_),
    .X(_00050_));
 a22o_1 _15575_ (.A1(net439),
    .A2(_07114_),
    .B1(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_key_o ),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[2] ),
    .X(_00049_));
 o211a_1 _15576_ (.A1(_10732_),
    .A2(_10734_),
    .B1(net473),
    .C1(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_3b_o ),
    .X(_10737_));
 and3_1 _15577_ (.A(net470),
    .B(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_2b_o ),
    .C(_10731_),
    .X(_10738_));
 a21o_1 _15578_ (.A1(net463),
    .A2(_07114_),
    .B1(_10738_),
    .X(_10739_));
 or2_1 _15579_ (.A(_10737_),
    .B(_10739_),
    .X(_00048_));
 nor2_1 _15580_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[0] ),
    .B(_07520_),
    .Y(_10740_));
 a21o_2 _15581_ (.A1(\digitop_pav2.sec_inst.ld_mem.st[2] ),
    .A2(net714),
    .B1(_07568_),
    .X(_10741_));
 a21o_1 _15582_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[2] ),
    .A2(_10741_),
    .B1(_07517_),
    .X(_10742_));
 a311o_2 _15583_ (.A1(_07093_),
    .A2(_10421_),
    .A3(_10740_),
    .B1(_10742_),
    .C1(net463),
    .X(_10743_));
 inv_2 _15584_ (.A(_10743_),
    .Y(_10744_));
 a22o_1 _15585_ (.A1(net426),
    .A2(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_2b_o ),
    .B1(net413),
    .B2(net463),
    .X(_10745_));
 o21a_1 _15586_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[4] ),
    .A2(net439),
    .B1(net413),
    .X(_10746_));
 a211o_1 _15587_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_key_o ),
    .B1(_10745_),
    .C1(_10746_),
    .X(_10747_));
 or2_1 _15588_ (.A(net373),
    .B(_10747_),
    .X(_10748_));
 o32a_1 _15589_ (.A1(_10737_),
    .A2(_10738_),
    .A3(_10748_),
    .B1(_10421_),
    .B2(net366),
    .X(_10749_));
 inv_2 _15590_ (.A(_10749_),
    .Y(_10750_));
 or2_1 _15591_ (.A(_10743_),
    .B(_10749_),
    .X(_10751_));
 o31ai_1 _15592_ (.A1(_07518_),
    .A2(_10421_),
    .A3(_10751_),
    .B1(net413),
    .Y(_10752_));
 a22o_1 _15593_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[0] ),
    .A2(_10421_),
    .B1(_10752_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[4] ),
    .X(_00047_));
 and3_1 _15594_ (.A(net463),
    .B(_10732_),
    .C(_10735_),
    .X(_10753_));
 and4_1 _15595_ (.A(net473),
    .B(net413),
    .C(_10731_),
    .D(_10735_),
    .X(_10754_));
 and2_1 _15596_ (.A(net470),
    .B(_07112_),
    .X(_10755_));
 a211o_1 _15597_ (.A1(net413),
    .A2(_10753_),
    .B1(_10754_),
    .C1(_10755_),
    .X(_00046_));
 a2bb2o_1 _15598_ (.A1_N(_07093_),
    .A2_N(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_key_o ),
    .B1(net413),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[4] ),
    .X(_00045_));
 mux2_1 _15599_ (.A0(net473),
    .A1(net439),
    .S(net413),
    .X(_10756_));
 a31o_1 _15600_ (.A1(net426),
    .A2(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_2b_o ),
    .A3(_10422_),
    .B1(_10756_),
    .X(_00044_));
 or2_1 _15601_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[4] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[6] ),
    .X(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_form_enable ));
 and3_1 _15602_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[0] ),
    .B(net159),
    .C(_07846_),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_rd_stb ));
 or2_1 _15603_ (.A(_09501_),
    .B(\digitop_pav2.testctrl_pav2.inst_mode.n_state[0] ),
    .X(_10757_));
 nor2_1 _15604_ (.A(_09492_),
    .B(_10757_),
    .Y(_10758_));
 and3_1 _15605_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.n_state[4] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mode.n_state[2] ),
    .C(_10758_),
    .X(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_mbist ));
 nand2_1 _15606_ (.A(net1309),
    .B(\digitop_pav2.testctrl_pav2.inst_mode.n_state[0] ),
    .Y(_10759_));
 nor2_1 _15607_ (.A(_09491_),
    .B(_10759_),
    .Y(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_dummy ));
 or2_1 _15608_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.n_state[1] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mode.n_state[0] ),
    .X(_10760_));
 nor2_1 _15609_ (.A(_09491_),
    .B(_10760_),
    .Y(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_probe ));
 or3b_1 _15610_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.n_state[2] ),
    .B(_09501_),
    .C_N(\digitop_pav2.testctrl_pav2.inst_mode.n_state[0] ),
    .X(_10761_));
 nand2_1 _15611_ (.A(_09459_),
    .B(_09492_),
    .Y(_10762_));
 nor2_1 _15612_ (.A(_10761_),
    .B(_10762_),
    .Y(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_anafunc ));
 or2_1 _15613_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.n_state[2] ),
    .B(_10762_),
    .X(_10763_));
 nor2_1 _15614_ (.A(_10757_),
    .B(_10763_),
    .Y(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_digfunc ));
 nor2_1 _15615_ (.A(_10759_),
    .B(_10763_),
    .Y(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_calclk ));
 nand2_1 _15616_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.n_state[2] ),
    .B(_09492_),
    .Y(_10764_));
 a21bo_1 _15617_ (.A1(\digitop_pav2.testctrl_pav2.inst_mode.n_state[2] ),
    .A2(net1309),
    .B1_N(_10761_),
    .X(_10765_));
 o2bb2a_1 _15618_ (.A1_N(\digitop_pav2.testctrl_pav2.inst_mode.n_state[3] ),
    .A2_N(_10765_),
    .B1(_10764_),
    .B2(_10757_),
    .X(_10766_));
 nor2_1 _15619_ (.A(_09459_),
    .B(_10766_),
    .Y(_10767_));
 or4_1 _15620_ (.A(_09480_),
    .B(_09486_),
    .C(_09511_),
    .D(_10767_),
    .X(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_clkout ));
 o31a_1 _15621_ (.A1(_07084_),
    .A2(net1486),
    .A3(_09453_),
    .B1(_09494_),
    .X(_10768_));
 o211ai_1 _15622_ (.A1(_09491_),
    .A2(_10757_),
    .B1(_10768_),
    .C1(_09426_),
    .Y(_10769_));
 a31o_1 _15623_ (.A1(\digitop_pav2.testctrl_pav2.inst_mode.n_state[4] ),
    .A2(_09492_),
    .A3(_10765_),
    .B1(_10769_),
    .X(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_rnclkout ));
 and3_1 _15624_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.tm_amux ),
    .B(_09432_),
    .C(_09463_),
    .X(_00165_));
 and3_1 _15625_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.tm_amux ),
    .B(_09463_),
    .C(_09475_),
    .X(_00166_));
 and3_1 _15626_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.tm_amux ),
    .B(_09456_),
    .C(_09463_),
    .X(_00167_));
 and3_1 _15627_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.tm_amux ),
    .B(_09439_),
    .C(_09463_),
    .X(_00164_));
 and3_1 _15628_ (.A(_07084_),
    .B(_09430_),
    .C(_09439_),
    .X(_10770_));
 o21a_1 _15629_ (.A1(_09463_),
    .A2(_10770_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mode.tm_amux ),
    .X(_00163_));
 or3_1 _15630_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_state[2] ),
    .B(_00114_),
    .C(_00115_),
    .X(_10771_));
 nor2_1 _15631_ (.A(_00113_),
    .B(_10771_),
    .Y(_10772_));
 and2_1 _15632_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[4] ),
    .B(_10772_),
    .X(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_int_rd_end ));
 and2_1 _15633_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[1] ),
    .B(_10772_),
    .X(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_int_wr_end ));
 or2_2 _15634_ (.A(net1727),
    .B(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_9.Y ),
    .X(\digitop_pav2.pass_t2 ));
 and3_2 _15635_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_mode_after_buf ),
    .B(net192),
    .C(net530),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.int_rst_b ));
 and3b_1 _15636_ (.A_N(\digitop_pav2.sync_inst.inst_clkx.inst_cipher.inst_en.cipher_off_ff ),
    .B(net1244),
    .C(_09160_),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cipher.cipher_en ));
 or4_1 _15637_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[3] ),
    .B(net464),
    .C(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_key_o ),
    .D(_07517_),
    .X(_10773_));
 a21o_1 _15638_ (.A1(net426),
    .A2(_10422_),
    .B1(_10773_),
    .X(_00130_));
 a2111o_1 _15639_ (.A1(net464),
    .A2(net413),
    .B1(_10755_),
    .C1(_10756_),
    .D1(net426),
    .X(_10774_));
 a21oi_1 _15640_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[3] ),
    .A2(_10732_),
    .B1(_10774_),
    .Y(_10775_));
 xnor2_1 _15641_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[2] ),
    .B(_08909_),
    .Y(_10776_));
 a2bb2o_1 _15642_ (.A1_N(_10775_),
    .A2_N(_10776_),
    .B1(_08880_),
    .B2(_00049_),
    .X(_10777_));
 xnor2_1 _15643_ (.A(_07106_),
    .B(_10777_),
    .Y(_10778_));
 xnor2_1 _15644_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[1] ),
    .B(_08913_),
    .Y(_10779_));
 o2bb2a_1 _15645_ (.A1_N(_08881_),
    .A2_N(_00049_),
    .B1(_10775_),
    .B2(_10779_),
    .X(_10780_));
 nor2_1 _15646_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[1] ),
    .B(_10780_),
    .Y(_10781_));
 xnor2_1 _15647_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[0] ),
    .B(_08908_),
    .Y(_10782_));
 a2bb2o_1 _15648_ (.A1_N(_10775_),
    .A2_N(_10782_),
    .B1(_08883_),
    .B2(_00049_),
    .X(_10783_));
 and2_1 _15649_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[1] ),
    .B(_10780_),
    .X(_10784_));
 mux2_1 _15650_ (.A0(_10781_),
    .A1(_10784_),
    .S(_10778_),
    .X(_10785_));
 nor2_1 _15651_ (.A(_10744_),
    .B(_10749_),
    .Y(_10786_));
 xor2_1 _15652_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[0] ),
    .B(_10783_),
    .X(_10787_));
 o31ai_1 _15653_ (.A1(_10778_),
    .A2(_10781_),
    .A3(_10784_),
    .B1(_10783_),
    .Y(_10788_));
 o2111a_1 _15654_ (.A1(_10783_),
    .A2(_10785_),
    .B1(_10786_),
    .C1(_10787_),
    .D1(_10788_),
    .X(_00128_));
 nor4_1 _15655_ (.A(net473),
    .B(_10739_),
    .C(_10753_),
    .D(_10755_),
    .Y(_10789_));
 nor3_2 _15656_ (.A(net427),
    .B(_10733_),
    .C(_10736_),
    .Y(_10790_));
 o221a_1 _15657_ (.A1(_08911_),
    .A2(_10789_),
    .B1(_10790_),
    .B2(_08897_),
    .C1(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[1] ),
    .X(_10791_));
 o221a_1 _15658_ (.A1(_08912_),
    .A2(net335),
    .B1(_10790_),
    .B2(_08898_),
    .C1(_07040_),
    .X(_10792_));
 nor2_1 _15659_ (.A(_10791_),
    .B(_10792_),
    .Y(_10793_));
 xnor2_1 _15660_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_0.A ),
    .B(_10793_),
    .Y(_10794_));
 o22a_1 _15661_ (.A1(_08903_),
    .A2(net335),
    .B1(_10790_),
    .B2(_08900_),
    .X(_10795_));
 o22a_1 _15662_ (.A1(_08904_),
    .A2(net335),
    .B1(_10790_),
    .B2(_08901_),
    .X(_10796_));
 mux2_1 _15663_ (.A0(_10796_),
    .A1(_10795_),
    .S(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[0] ),
    .X(_10797_));
 or2_1 _15664_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_0.A ),
    .B(_10797_),
    .X(_10798_));
 or3_2 _15665_ (.A(_10733_),
    .B(_10745_),
    .C(_10754_),
    .X(_10799_));
 nand2_1 _15666_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_0.A ),
    .B(_10797_),
    .Y(_10800_));
 mux2_1 _15667_ (.A0(_10798_),
    .A1(_10800_),
    .S(_10794_),
    .X(_10801_));
 nor2_1 _15668_ (.A(_10799_),
    .B(_10801_),
    .Y(_00129_));
 and4bb_1 _15669_ (.A_N(_10794_),
    .B_N(_10799_),
    .C(_10800_),
    .D(_10798_),
    .X(_00126_));
 and3b_1 _15670_ (.A_N(_10787_),
    .B(_10786_),
    .C(_10785_),
    .X(_00127_));
 and2b_1 _15671_ (.A_N(ff_erase_ff3),
    .B(ff_erase_ff2),
    .X(ff_erase_rise));
 and2b_1 _15672_ (.A_N(ff_prog_ff3),
    .B(ff_prog_ff2),
    .X(ff_prog_rise));
 nor2_1 _15673_ (.A(net1481),
    .B(\digitop_pav2.testctrl_pav2.inst_mode.tm_digfunc ),
    .Y(_10802_));
 mux2_1 _15674_ (.A0(tclk_i),
    .A1(clk_i),
    .S(_10802_),
    .X(\digitop_pav2.func_clk_pre ));
 or4_1 _15675_ (.A(net1483),
    .B(\digitop_pav2.testctrl_pav2.inst_mode.tm_anafunc ),
    .C(\digitop_pav2.testctrl_pav2.inst_mode.tm_probe ),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.tm_dummy ),
    .X(_10803_));
 or4_1 _15676_ (.A(net1481),
    .B(\digitop_pav2.testctrl_pav2.inst_mode.tm_digfunc ),
    .C(\digitop_pav2.testctrl_pav2.inst_mode.tm_rnclkout ),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.tm_clkout ),
    .X(_10804_));
 a211oi_2 _15677_ (.A1(\digitop_pav2.testctrl_pav2.inst_enter.tm_enter ),
    .A2(_07163_),
    .B1(_10803_),
    .C1(_10804_),
    .Y(net140));
 mux2_1 _15678_ (.A0(clk_i),
    .A1(rnclk_i),
    .S(\digitop_pav2.testctrl_pav2.inst_mode.tm_rnclkout ),
    .X(_10805_));
 o21a_2 _15679_ (.A1(\digitop_pav2.testctrl_pav2.inst_mode.tm_rnclkout ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mode.tm_clkout ),
    .B1(_10805_),
    .X(_10806_));
 a211oi_1 _15680_ (.A1(net1481),
    .A2(_07169_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mode.tm_clkout ),
    .C1(\digitop_pav2.testctrl_pav2.inst_mode.tm_rnclkout ),
    .Y(_10807_));
 a21o_2 _15681_ (.A1(\digitop_pav2.fm0miller_inst.fm0x_mask.gand_delay ),
    .A2(\digitop_pav2.fm0miller_inst.fm0x_mask.tx_raw_i ),
    .B1(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[9].fm0miller_pav2_gor_dly.Y ),
    .X(_10808_));
 nand2_1 _15682_ (.A(net192),
    .B(_07167_),
    .Y(net78));
 o22a_2 _15683_ (.A1(net192),
    .A2(net1),
    .B1(_10808_),
    .B2(net78),
    .X(_10809_));
 o32a_2 _15684_ (.A1(net1481),
    .A2(_07168_),
    .A3(_10809_),
    .B1(_10807_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mode.tm_anafunc ),
    .X(_10810_));
 o22a_2 _15685_ (.A1(_07167_),
    .A2(net1),
    .B1(_10806_),
    .B2(_10810_),
    .X(_10811_));
 mux2_1 _15686_ (.A0(_10808_),
    .A1(_10811_),
    .S(_07113_),
    .X(_10812_));
 mux2_1 _15687_ (.A0(_10812_),
    .A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.calx_end_o ),
    .S(net1483),
    .X(net141));
 nand2_2 _15688_ (.A(net1481),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[2] ),
    .Y(_10813_));
 mux2_1 _15689_ (.A0(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[1] ),
    .A1(\digitop_pav2.memctrl_inst.bit_addr[1] ),
    .S(_10813_),
    .X(_10814_));
 mux2_2 _15690_ (.A0(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[0] ),
    .A1(\digitop_pav2.memctrl_inst.bit_addr[0] ),
    .S(_10813_),
    .X(_10815_));
 inv_2 _15691_ (.A(_10815_),
    .Y(_10816_));
 nor2_1 _15692_ (.A(net1024),
    .B(_10815_),
    .Y(_10817_));
 mux2_2 _15693_ (.A0(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[2] ),
    .A1(\digitop_pav2.memctrl_inst.bit_addr[2] ),
    .S(_10813_),
    .X(_10818_));
 or3_1 _15694_ (.A(net1024),
    .B(_10815_),
    .C(net1023),
    .X(_10819_));
 a21boi_1 _15695_ (.A1(\digitop_pav2.memctrl_inst.bit_addr_allow ),
    .A2(_09383_),
    .B1_N(_10813_),
    .Y(_10820_));
 a21bo_1 _15696_ (.A1(\digitop_pav2.memctrl_inst.bit_addr_allow ),
    .A2(_09383_),
    .B1_N(_10813_),
    .X(_10821_));
 mux2_2 _15697_ (.A0(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[3] ),
    .A1(\digitop_pav2.memctrl_inst.bit_addr[3] ),
    .S(_10813_),
    .X(_10822_));
 nor2_2 _15698_ (.A(_10820_),
    .B(_10822_),
    .Y(_10823_));
 or2_2 _15699_ (.A(_10820_),
    .B(_10822_),
    .X(_10824_));
 nor2_1 _15700_ (.A(_10819_),
    .B(_10824_),
    .Y(net88));
 or3_1 _15701_ (.A(net1024),
    .B(_10816_),
    .C(net1023),
    .X(_10825_));
 or2_2 _15702_ (.A(_10824_),
    .B(_10825_),
    .X(_10826_));
 inv_2 _15703_ (.A(_10826_),
    .Y(net95));
 or3b_1 _15704_ (.A(net1023),
    .B(_10815_),
    .C_N(net1024),
    .X(_10827_));
 nor2_2 _15705_ (.A(_10824_),
    .B(_10827_),
    .Y(net96));
 and3b_1 _15706_ (.A_N(net1023),
    .B(net1024),
    .C(_10815_),
    .X(_10828_));
 nand2_2 _15707_ (.A(_10823_),
    .B(_10828_),
    .Y(_10829_));
 inv_2 _15708_ (.A(_10829_),
    .Y(net97));
 and3_2 _15709_ (.A(_10817_),
    .B(net1023),
    .C(_10823_),
    .X(net98));
 or4b_4 _15710_ (.A(_10814_),
    .B(_10824_),
    .C(_10816_),
    .D_N(net1023),
    .X(_10830_));
 inv_2 _15711_ (.A(_10830_),
    .Y(net99));
 and4_2 _15712_ (.A(net1024),
    .B(_10816_),
    .C(net1023),
    .D(_10823_),
    .X(net100));
 and4_1 _15713_ (.A(net1024),
    .B(_10815_),
    .C(net1023),
    .D(_10823_),
    .X(net101));
 and2_2 _15714_ (.A(_10821_),
    .B(_10822_),
    .X(_10831_));
 nand2_2 _15715_ (.A(_10821_),
    .B(_10822_),
    .Y(_10832_));
 or2_2 _15716_ (.A(_10819_),
    .B(_10832_),
    .X(_10833_));
 inv_2 _15717_ (.A(_10833_),
    .Y(net102));
 or2_1 _15718_ (.A(_10825_),
    .B(_10832_),
    .X(_10834_));
 inv_2 _15719_ (.A(_10834_),
    .Y(net103));
 nor2_2 _15720_ (.A(_10827_),
    .B(_10832_),
    .Y(net89));
 nand2_4 _15721_ (.A(_10828_),
    .B(_10831_),
    .Y(_10835_));
 inv_2 _15722_ (.A(_10835_),
    .Y(net90));
 and3_2 _15723_ (.A(_10817_),
    .B(net1023),
    .C(_10831_),
    .X(net91));
 or4b_2 _15724_ (.A(net1024),
    .B(_10832_),
    .C(_10816_),
    .D_N(net1023),
    .X(_10836_));
 inv_2 _15725_ (.A(_10836_),
    .Y(net92));
 and4_2 _15726_ (.A(net1024),
    .B(_10816_),
    .C(_10818_),
    .D(_10831_),
    .X(net93));
 and4_2 _15727_ (.A(net1024),
    .B(_10815_),
    .C(_10818_),
    .D(_10831_),
    .X(net94));
 o21a_1 _15728_ (.A1(net1491),
    .A2(_09450_),
    .B1(_09476_),
    .X(_10837_));
 mux2_2 _15729_ (.A0(_07097_),
    .A1(\digitop_pav2.cal_inst.calx_mux.dtest_trim_0_i ),
    .S(net1482),
    .X(_10838_));
 mux2_1 _15730_ (.A0(_10838_),
    .A1(_10837_),
    .S(\digitop_pav2.testctrl_pav2.inst_mode.tm_clkout ),
    .X(net75));
 mux2_2 _15731_ (.A0(_07098_),
    .A1(\digitop_pav2.cal_inst.calx_mux.dtest_trim_1_i ),
    .S(net1482),
    .X(_10839_));
 mux2_1 _15732_ (.A0(_10839_),
    .A1(_09431_),
    .S(\digitop_pav2.testctrl_pav2.inst_mode.tm_clkout ),
    .X(net76));
 mux2_2 _15733_ (.A0(\digitop_pav2.access_inst.access_check0.fg_i[7] ),
    .A1(\digitop_pav2.cal_inst.calx_mux.dtest_trim_2_i ),
    .S(net1482),
    .X(_10840_));
 mux2_1 _15734_ (.A0(_10840_),
    .A1(_09454_),
    .S(\digitop_pav2.testctrl_pav2.inst_mode.tm_clkout ),
    .X(net77));
 o21a_1 _15735_ (.A1(net1491),
    .A2(_09426_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mode.tm_rnclkout ),
    .X(_10841_));
 a2bb2o_1 _15736_ (.A1_N(net1324),
    .A2_N(\digitop_pav2.testctrl_pav2.inst_mode.tm_rnclkout ),
    .B1(_09508_),
    .B2(_10841_),
    .X(net81));
 mux2_1 _15737_ (.A0(_07095_),
    .A1(_09428_),
    .S(\digitop_pav2.testctrl_pav2.inst_mode.tm_rnclkout ),
    .X(net82));
 and2b_1 _15738_ (.A_N(\digitop_pav2.testctrl_pav2.inst_mode.tm_rnclkout ),
    .B(\digitop_pav2.access_inst.access_check0.fg_i[2] ),
    .X(_10842_));
 a41o_1 _15739_ (.A1(\digitop_pav2.testctrl_pav2.inst_mode.tm_rnclkout ),
    .A2(_09424_),
    .A3(_09442_),
    .A4(_09453_),
    .B1(_10842_),
    .X(net83));
 or2_1 _15740_ (.A(net1503),
    .B(_07167_),
    .X(_10843_));
 o211a_2 _15741_ (.A1(\digitop_pav2.testctrl_pav2.inst_mode.tm_anafunc ),
    .A2(_10808_),
    .B1(_10843_),
    .C1(_07113_),
    .X(net79));
 and3_2 _15742_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_mode_after_buf ),
    .B(net192),
    .C(_09538_),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.cp_div_sel[0] ));
 and3_2 _15743_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_mode_after_buf ),
    .B(net192),
    .C(_09537_),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.cp_div_sel[1] ));
 mux2_1 _15744_ (.A0(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.scwend_clk_i ),
    .A1(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.boot_dis_clk_after_buf ),
    .S(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.en_pup_clk_b ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_trigger.trigger_clk ));
 and3_1 _15745_ (.A(_07130_),
    .B(_07170_),
    .C(\digitop_pav2.proc_ctrl_inst.int_pass_t2_flag ),
    .X(_00145_));
 and2b_1 _15746_ (.A_N(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_9.Y ),
    .B(_09087_),
    .X(_00144_));
 and3_1 _15747_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[0] ),
    .B(net426),
    .C(\digitop_pav2.aes128_inst.aes128_counter.cnt_rnd_en_o ),
    .X(_10844_));
 a21o_1 _15748_ (.A1(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[1] ),
    .A2(_10844_),
    .B1(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[2] ),
    .X(_10845_));
 and3_1 _15749_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[1] ),
    .C(_10844_),
    .X(_10846_));
 or3b_2 _15750_ (.A(_10846_),
    .B(_10741_),
    .C_N(_10845_),
    .X(_10847_));
 inv_2 _15751_ (.A(_10847_),
    .Y(_01286_));
 a21oi_1 _15752_ (.A1(net426),
    .A2(\digitop_pav2.aes128_inst.aes128_counter.cnt_rnd_en_o ),
    .B1(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[0] ),
    .Y(_10848_));
 nor3_2 _15753_ (.A(_10741_),
    .B(_10844_),
    .C(_10848_),
    .Y(_01284_));
 xnor2_1 _15754_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[1] ),
    .B(_10844_),
    .Y(_10849_));
 nor2_1 _15755_ (.A(_10741_),
    .B(_10849_),
    .Y(_01285_));
 nor2_1 _15756_ (.A(_01284_),
    .B(_01285_),
    .Y(_10850_));
 and2_1 _15757_ (.A(_10847_),
    .B(_10850_),
    .X(_00000_));
 or3b_1 _15758_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[1] ),
    .B(_01286_),
    .C_N(_01284_),
    .X(_10851_));
 inv_2 _15759_ (.A(_10851_),
    .Y(_10852_));
 o21bai_1 _15760_ (.A1(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[3] ),
    .A2(_10846_),
    .B1_N(_10741_),
    .Y(_10853_));
 a21oi_2 _15761_ (.A1(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[3] ),
    .A2(_10846_),
    .B1(_10853_),
    .Y(_01287_));
 a31o_1 _15762_ (.A1(_10847_),
    .A2(_10849_),
    .A3(_01287_),
    .B1(_10852_),
    .X(_00001_));
 and2_1 _15763_ (.A(_10852_),
    .B(_01287_),
    .X(_10854_));
 and2b_1 _15764_ (.A_N(_01284_),
    .B(_01285_),
    .X(_10855_));
 nor2_1 _15765_ (.A(_01286_),
    .B(_01287_),
    .Y(_10856_));
 a21o_1 _15766_ (.A1(_10855_),
    .A2(_10856_),
    .B1(_10854_),
    .X(_00002_));
 a32o_1 _15767_ (.A1(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[1] ),
    .A2(_01284_),
    .A3(_10856_),
    .B1(_01287_),
    .B2(_00000_),
    .X(_00003_));
 nor2_1 _15768_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[3] ),
    .B(_10847_),
    .Y(_10857_));
 a32o_1 _15769_ (.A1(_10847_),
    .A2(_10849_),
    .A3(_01287_),
    .B1(_10857_),
    .B2(_10850_),
    .X(_00004_));
 a31o_1 _15770_ (.A1(_07040_),
    .A2(_01284_),
    .A3(_10857_),
    .B1(_10854_),
    .X(_00005_));
 o31a_1 _15771_ (.A1(net188),
    .A2(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[3] ),
    .A3(_09563_),
    .B1(_09552_),
    .X(_10858_));
 or3b_1 _15772_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[3] ),
    .B(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[2] ),
    .C_N(_09553_),
    .X(_10859_));
 a31o_1 _15773_ (.A1(net188),
    .A2(_09551_),
    .A3(_10859_),
    .B1(_10858_),
    .X(_10860_));
 inv_2 _15774_ (.A(_10860_),
    .Y(_10861_));
 nand2_1 _15775_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[3] ),
    .B(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[2] ),
    .Y(_10862_));
 and2_1 _15776_ (.A(_09552_),
    .B(_10859_),
    .X(_10863_));
 a31o_1 _15777_ (.A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[3] ),
    .A2(_09551_),
    .A3(_09563_),
    .B1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[4] ),
    .X(_10864_));
 o22a_1 _15778_ (.A1(_08520_),
    .A2(_10861_),
    .B1(_10863_),
    .B2(_10864_),
    .X(_10865_));
 and4b_1 _15779_ (.A_N(_09563_),
    .B(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[4] ),
    .C(_09551_),
    .D(_10859_),
    .X(_10866_));
 a41o_1 _15780_ (.A1(_07122_),
    .A2(_09561_),
    .A3(_10858_),
    .A4(_10862_),
    .B1(net531),
    .X(_10867_));
 a221o_1 _15781_ (.A1(_08520_),
    .A2(_10860_),
    .B1(_10866_),
    .B2(_07124_),
    .C1(_10867_),
    .X(_10868_));
 o21a_1 _15782_ (.A1(net530),
    .A2(_10865_),
    .B1(_10868_),
    .X(\digitop_pav2.fm0miller_inst.fm0x_ctrl.n_dt_tx_st ));
 and2_1 _15783_ (.A(net191),
    .B(net192),
    .X(\digitop_pav2.fm0miller_inst.ctrl[0] ));
 and2_1 _15784_ (.A(net190),
    .B(net192),
    .X(\digitop_pav2.fm0miller_inst.ctrl[1] ));
 and2_1 _15785_ (.A(net189),
    .B(net192),
    .X(\digitop_pav2.fm0miller_inst.ctrl[2] ));
 nor2_1 _15786_ (.A(_07244_),
    .B(_07275_),
    .Y(_10869_));
 o22a_1 _15787_ (.A1(_07244_),
    .A2(_07275_),
    .B1(_08488_),
    .B2(_07274_),
    .X(_10870_));
 a22o_1 _15788_ (.A1(_07257_),
    .A2(_07363_),
    .B1(_10870_),
    .B2(_07278_),
    .X(_10871_));
 and2b_1 _15789_ (.A_N(_10460_),
    .B(_10871_),
    .X(_10872_));
 a32o_1 _15790_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[5] ),
    .A2(_07330_),
    .A3(_10498_),
    .B1(net1162),
    .B2(net1289),
    .X(_10873_));
 or2_1 _15791_ (.A(_10499_),
    .B(_10873_),
    .X(_10874_));
 o221a_1 _15792_ (.A1(_07347_),
    .A2(net1229),
    .B1(_10480_),
    .B2(_10514_),
    .C1(_07293_),
    .X(_10875_));
 or4_1 _15793_ (.A(_10525_),
    .B(_10872_),
    .C(_10874_),
    .D(_10875_),
    .X(\digitop_pav2.proc_ctrl_inst.cmdfsm.n_rn_rst_b ));
 a21oi_1 _15794_ (.A1(_07244_),
    .A2(_08488_),
    .B1(_07279_),
    .Y(_10876_));
 a31o_1 _15795_ (.A1(_07274_),
    .A2(_10530_),
    .A3(_10876_),
    .B1(_10515_),
    .X(\digitop_pav2.proc_ctrl_inst.cmdfsm.n_rn_en ));
 nand2_1 _15796_ (.A(net1241),
    .B(_09096_),
    .Y(_10877_));
 and2_2 _15797_ (.A(_07160_),
    .B(_09146_),
    .X(_10878_));
 nand2_4 _15798_ (.A(_07160_),
    .B(_09146_),
    .Y(_10879_));
 nor2_1 _15799_ (.A(net1233),
    .B(_10879_),
    .Y(_10880_));
 nand2_1 _15800_ (.A(net1245),
    .B(_10878_),
    .Y(_10881_));
 a31o_1 _15801_ (.A1(net1246),
    .A2(_07160_),
    .A3(_09144_),
    .B1(_10877_),
    .X(_10882_));
 nor2_1 _15802_ (.A(net1241),
    .B(_09097_),
    .Y(_10883_));
 or2_2 _15803_ (.A(net1241),
    .B(_09097_),
    .X(_10884_));
 o21a_1 _15804_ (.A1(_10880_),
    .A2(_10884_),
    .B1(_10882_),
    .X(_10885_));
 nor2_1 _15805_ (.A(\digitop_pav2.proc_ctrl_inst.profsm.r1_ff ),
    .B(_08870_),
    .Y(_10886_));
 a21oi_1 _15806_ (.A1(_07243_),
    .A2(net1225),
    .B1(net1246),
    .Y(_10887_));
 nor2_1 _15807_ (.A(net969),
    .B(_07244_),
    .Y(_10888_));
 a211o_1 _15808_ (.A1(net969),
    .A2(_10692_),
    .B1(_10888_),
    .C1(net1246),
    .X(_10889_));
 o41a_1 _15809_ (.A1(net1233),
    .A2(net968),
    .A3(net1163),
    .A4(_10886_),
    .B1(_10889_),
    .X(_10890_));
 a2bb2o_1 _15810_ (.A1_N(_10885_),
    .A2_N(_10890_),
    .B1(net1187),
    .B2(_09096_),
    .X(_10891_));
 and2_1 _15811_ (.A(_09031_),
    .B(_10693_),
    .X(_10892_));
 or4b_1 _15812_ (.A(net1247),
    .B(net969),
    .C(\digitop_pav2.proc_ctrl_inst.profsm.skip_abort ),
    .D_N(\digitop_pav2.proc_ctrl_inst.int_pass_t2_flag ),
    .X(_10893_));
 nand2_1 _15813_ (.A(_10892_),
    .B(_10893_),
    .Y(_10894_));
 o21a_1 _15814_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.pro_abort_b_i ),
    .A2(_10692_),
    .B1(_10894_),
    .X(_10895_));
 nor2_1 _15815_ (.A(net1186),
    .B(_10879_),
    .Y(_10896_));
 or3b_1 _15816_ (.A(\digitop_pav2.proc_ctrl_inst.int_pass_t2_flag ),
    .B(_07311_),
    .C_N(_09149_),
    .X(_10897_));
 a32o_1 _15817_ (.A1(_09151_),
    .A2(_10879_),
    .A3(_10897_),
    .B1(_10896_),
    .B2(_10698_),
    .X(_10898_));
 and3_1 _15818_ (.A(net1246),
    .B(\digitop_pav2.proc_ctrl_inst.cmdctr.pro_abort_b_i ),
    .C(_10898_),
    .X(_10899_));
 o221a_1 _15819_ (.A1(_07130_),
    .A2(net969),
    .B1(_10895_),
    .B2(_10899_),
    .C1(_10695_),
    .X(_10900_));
 o22a_1 _15820_ (.A1(net969),
    .A2(_09031_),
    .B1(_10891_),
    .B2(_10900_),
    .X(_10901_));
 nor2_1 _15821_ (.A(net1246),
    .B(net968),
    .Y(_10902_));
 or2_1 _15822_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[1] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[2] ),
    .X(_10903_));
 or3b_1 _15823_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[1] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[2] ),
    .C_N(net1241),
    .X(_10904_));
 a21o_1 _15824_ (.A1(net1163),
    .A2(_10879_),
    .B1(net1233),
    .X(_10905_));
 o21ai_2 _15825_ (.A1(net1233),
    .A2(net968),
    .B1(_10905_),
    .Y(_10906_));
 o31a_1 _15826_ (.A1(net968),
    .A2(net1163),
    .A3(_10878_),
    .B1(_10906_),
    .X(_10907_));
 o21a_1 _15827_ (.A1(_07292_),
    .A2(_09149_),
    .B1(_09147_),
    .X(_10908_));
 and2_1 _15828_ (.A(_10879_),
    .B(_10908_),
    .X(_10909_));
 xnor2_1 _15829_ (.A(net969),
    .B(_10909_),
    .Y(_10910_));
 or2_4 _15830_ (.A(net1241),
    .B(_10903_),
    .X(_10911_));
 inv_2 _15831_ (.A(_10911_),
    .Y(_10912_));
 a2bb2o_1 _15832_ (.A1_N(net1196),
    .A2_N(_10881_),
    .B1(_10910_),
    .B2(net1244),
    .X(_10913_));
 o22a_1 _15833_ (.A1(_10904_),
    .A2(_10907_),
    .B1(_10911_),
    .B2(_10913_),
    .X(_10914_));
 nor2_1 _15834_ (.A(_10902_),
    .B(_10914_),
    .Y(_10915_));
 a311o_1 _15835_ (.A1(\digitop_pav2.proc_ctrl_inst.int_timeout_t2 ),
    .A2(\digitop_pav2.proc_ctrl_inst.cmdctr.pro_abort_b_i ),
    .A3(_10695_),
    .B1(_10901_),
    .C1(_10915_),
    .X(\digitop_pav2.proc_ctrl_inst.profsm.n_blf_abort ));
 nand2_1 _15836_ (.A(\digitop_pav2.pie_inst.fsm.temptari[9] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[6] ),
    .Y(_10916_));
 inv_2 _15837_ (.A(_10916_),
    .Y(_10917_));
 or2_1 _15838_ (.A(\digitop_pav2.pie_inst.fsm.temptari[9] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[6] ),
    .X(_10918_));
 nand2_1 _15839_ (.A(_10916_),
    .B(_10918_),
    .Y(_10919_));
 nand2_1 _15840_ (.A(\digitop_pav2.pie_inst.fsm.temptari[8] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[5] ),
    .Y(_10920_));
 or2_1 _15841_ (.A(\digitop_pav2.pie_inst.fsm.temptari[8] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[5] ),
    .X(_10921_));
 nand2_1 _15842_ (.A(_10920_),
    .B(_10921_),
    .Y(_10922_));
 nand2_1 _15843_ (.A(\digitop_pav2.pie_inst.fsm.temptari[7] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[4] ),
    .Y(_10923_));
 or2_1 _15844_ (.A(\digitop_pav2.pie_inst.fsm.temptari[7] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[4] ),
    .X(_10924_));
 nand2_1 _15845_ (.A(_10923_),
    .B(_10924_),
    .Y(_10925_));
 nand2_1 _15846_ (.A(\digitop_pav2.pie_inst.fsm.temptari[6] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[3] ),
    .Y(_10926_));
 or2_1 _15847_ (.A(\digitop_pav2.pie_inst.fsm.temptari[6] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[3] ),
    .X(_10927_));
 nand2_1 _15848_ (.A(_10926_),
    .B(_10927_),
    .Y(_10928_));
 nand2_1 _15849_ (.A(\digitop_pav2.pie_inst.fsm.temptari[5] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[2] ),
    .Y(_10929_));
 or2_1 _15850_ (.A(\digitop_pav2.pie_inst.fsm.temptari[5] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[2] ),
    .X(_10930_));
 nand2_1 _15851_ (.A(_10929_),
    .B(_10930_),
    .Y(_10931_));
 xor2_1 _15852_ (.A(\digitop_pav2.pie_inst.fsm.temptari[4] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[1] ),
    .X(_10932_));
 nand2_1 _15853_ (.A(\digitop_pav2.pie_inst.fsm.temptari[3] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[0] ),
    .Y(_10933_));
 and3_1 _15854_ (.A(\digitop_pav2.pie_inst.fsm.temptari[3] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[0] ),
    .C(_10932_),
    .X(_10934_));
 a21o_1 _15855_ (.A1(\digitop_pav2.pie_inst.fsm.temptari[4] ),
    .A2(\digitop_pav2.pie_inst.fsm.temptari[1] ),
    .B1(_10934_),
    .X(_10935_));
 a21bo_1 _15856_ (.A1(_10930_),
    .A2(_10935_),
    .B1_N(_10929_),
    .X(_10936_));
 a21boi_1 _15857_ (.A1(_10927_),
    .A2(_10936_),
    .B1_N(_10926_),
    .Y(_10937_));
 o21ai_1 _15858_ (.A1(_10925_),
    .A2(_10937_),
    .B1(_10923_),
    .Y(_10938_));
 a21boi_1 _15859_ (.A1(_10921_),
    .A2(_10938_),
    .B1_N(_10920_),
    .Y(_10939_));
 nor2_1 _15860_ (.A(_10919_),
    .B(_10939_),
    .Y(_10940_));
 o21a_1 _15861_ (.A1(_10917_),
    .A2(_10940_),
    .B1(\digitop_pav2.pie_inst.fsm.temptari[7] ),
    .X(_10941_));
 nor3_1 _15862_ (.A(\digitop_pav2.pie_inst.fsm.temptari[7] ),
    .B(_10917_),
    .C(_10940_),
    .Y(_10942_));
 nor2_1 _15863_ (.A(_10941_),
    .B(_10942_),
    .Y(_10943_));
 xor2_1 _15864_ (.A(_10919_),
    .B(_10939_),
    .X(_10944_));
 xor2_1 _15865_ (.A(_10922_),
    .B(_10938_),
    .X(_10945_));
 inv_2 _15866_ (.A(_10945_),
    .Y(_10946_));
 xor2_1 _15867_ (.A(_10925_),
    .B(_10937_),
    .X(_10947_));
 xor2_1 _15868_ (.A(_10928_),
    .B(_10936_),
    .X(_10948_));
 xnor2_4 _15869_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[4] ),
    .B(_09577_),
    .Y(_10949_));
 inv_2 _15870_ (.A(_10949_),
    .Y(\digitop_pav2.pie_inst.fsm.dif_pos_fix[4] ));
 xor2_1 _15871_ (.A(_10931_),
    .B(_10935_),
    .X(_10950_));
 and2b_1 _15872_ (.A_N(_10932_),
    .B(_10933_),
    .X(_10951_));
 nor2_1 _15873_ (.A(_10934_),
    .B(_10951_),
    .Y(_10952_));
 or2_1 _15874_ (.A(\digitop_pav2.pie_inst.fsm.temptari[3] ),
    .B(\digitop_pav2.pie_inst.fsm.temptari[0] ),
    .X(_10953_));
 and2_1 _15875_ (.A(_07146_),
    .B(\digitop_pav2.pie_inst.fsm.temptari[2] ),
    .X(_10954_));
 a22o_1 _15876_ (.A1(_10933_),
    .A2(_10953_),
    .B1(_10954_),
    .B2(_07147_),
    .X(_10955_));
 nand2_1 _15877_ (.A(\digitop_pav2.pie_inst.fsm.dif_pos_fix[0] ),
    .B(\digitop_pav2.pie_inst.fsm.past_ctr[1] ),
    .Y(_10956_));
 nand2_1 _15878_ (.A(_09573_),
    .B(_10956_),
    .Y(_10957_));
 inv_2 _15879_ (.A(_10957_),
    .Y(\digitop_pav2.pie_inst.fsm.dif_pos_fix[1] ));
 o221a_1 _15880_ (.A1(_09576_),
    .A2(_10952_),
    .B1(_10954_),
    .B2(_10957_),
    .C1(_10955_),
    .X(_10958_));
 a21oi_1 _15881_ (.A1(_09576_),
    .A2(_10952_),
    .B1(_10958_),
    .Y(_10959_));
 o21a_1 _15882_ (.A1(\digitop_pav2.pie_inst.fsm.dif_pos_fix[3] ),
    .A2(_10950_),
    .B1(_10959_),
    .X(_10960_));
 or2_1 _15883_ (.A(_10948_),
    .B(\digitop_pav2.pie_inst.fsm.dif_pos_fix[4] ),
    .X(_10961_));
 a221o_1 _15884_ (.A1(_10948_),
    .A2(\digitop_pav2.pie_inst.fsm.dif_pos_fix[4] ),
    .B1(_10950_),
    .B2(\digitop_pav2.pie_inst.fsm.dif_pos_fix[3] ),
    .C1(_10960_),
    .X(_10962_));
 o2bb2a_1 _15885_ (.A1_N(_10961_),
    .A2_N(_10962_),
    .B1(_09589_),
    .B2(_10947_),
    .X(_10963_));
 a221o_1 _15886_ (.A1(net493),
    .A2(_10946_),
    .B1(_10947_),
    .B2(_09589_),
    .C1(_10963_),
    .X(_10964_));
 o221a_1 _15887_ (.A1(_09581_),
    .A2(_10944_),
    .B1(_10946_),
    .B2(_09587_),
    .C1(_10964_),
    .X(_10965_));
 a221o_1 _15888_ (.A1(net491),
    .A2(_10943_),
    .B1(_10944_),
    .B2(net494),
    .C1(_10965_),
    .X(_10966_));
 or2_1 _15889_ (.A(\digitop_pav2.pie_inst.fsm.temptari[8] ),
    .B(_10941_),
    .X(_10967_));
 o221a_1 _15890_ (.A1(_09649_),
    .A2(_10943_),
    .B1(_10967_),
    .B2(_09585_),
    .C1(_10966_),
    .X(_10968_));
 a21bo_1 _15891_ (.A1(\digitop_pav2.pie_inst.fsm.past_ctr[2] ),
    .A2(\digitop_pav2.pie_inst.fsm.temptari[0] ),
    .B1_N(_09574_),
    .X(_10969_));
 a21o_1 _15892_ (.A1(\digitop_pav2.pie_inst.fsm.temptari[1] ),
    .A2(_10969_),
    .B1(_09583_),
    .X(_10970_));
 or2_1 _15893_ (.A(\digitop_pav2.pie_inst.fsm.temptari[1] ),
    .B(_10969_),
    .X(_10971_));
 a22o_1 _15894_ (.A1(\digitop_pav2.pie_inst.fsm.temptari[2] ),
    .A2(_10949_),
    .B1(_10970_),
    .B2(_10971_),
    .X(_10972_));
 o221a_1 _15895_ (.A1(\digitop_pav2.pie_inst.fsm.temptari[3] ),
    .A2(net495),
    .B1(_10949_),
    .B2(\digitop_pav2.pie_inst.fsm.temptari[2] ),
    .C1(_10972_),
    .X(_10973_));
 a221o_1 _15896_ (.A1(\digitop_pav2.pie_inst.fsm.temptari[4] ),
    .A2(net493),
    .B1(net495),
    .B2(\digitop_pav2.pie_inst.fsm.temptari[3] ),
    .C1(_10973_),
    .X(_10974_));
 o221a_1 _15897_ (.A1(\digitop_pav2.pie_inst.fsm.temptari[5] ),
    .A2(net494),
    .B1(_09587_),
    .B2(\digitop_pav2.pie_inst.fsm.temptari[4] ),
    .C1(_10974_),
    .X(_10975_));
 a221o_1 _15898_ (.A1(\digitop_pav2.pie_inst.fsm.temptari[5] ),
    .A2(net494),
    .B1(net491),
    .B2(\digitop_pav2.pie_inst.fsm.temptari[6] ),
    .C1(_10975_),
    .X(_10976_));
 o22a_1 _15899_ (.A1(\digitop_pav2.pie_inst.fsm.temptari[7] ),
    .A2(_09585_),
    .B1(net491),
    .B2(\digitop_pav2.pie_inst.fsm.temptari[6] ),
    .X(_10977_));
 a221o_1 _15900_ (.A1(\digitop_pav2.pie_inst.fsm.temptari[7] ),
    .A2(_09585_),
    .B1(_10976_),
    .B2(_10977_),
    .C1(\digitop_pav2.pie_inst.fsm.temptari[8] ),
    .X(_10978_));
 and4b_1 _15901_ (.A_N(\digitop_pav2.pie_inst.fsm.temptari[9] ),
    .B(\digitop_pav2.pie_inst.fsm.comp_delimiter_ff2 ),
    .C(_10978_),
    .D(\digitop_pav2.pie_inst.fsm.comp_tari_ff ),
    .X(_10979_));
 a21bo_1 _15902_ (.A1(\digitop_pav2.pie_inst.fsm.temptari[8] ),
    .A2(_10941_),
    .B1_N(_10979_),
    .X(_10980_));
 a211o_2 _15903_ (.A1(_09585_),
    .A2(_10967_),
    .B1(_10968_),
    .C1(_10980_),
    .X(_10981_));
 or2_1 _15904_ (.A(\digitop_pav2.pie_inst.fsm.pivot[2] ),
    .B(net495),
    .X(_10982_));
 o211a_1 _15905_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[1] ),
    .A2(_10949_),
    .B1(_09583_),
    .C1(\digitop_pav2.pie_inst.fsm.pivot[0] ),
    .X(_10983_));
 a221o_1 _15906_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[2] ),
    .A2(net495),
    .B1(_10949_),
    .B2(\digitop_pav2.pie_inst.fsm.pivot[1] ),
    .C1(_10983_),
    .X(_10984_));
 a22o_1 _15907_ (.A1(net1301),
    .A2(net493),
    .B1(_10982_),
    .B2(_10984_),
    .X(_10985_));
 o221a_1 _15908_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[4] ),
    .A2(net494),
    .B1(net493),
    .B2(net1301),
    .C1(_10985_),
    .X(_10986_));
 a221o_1 _15909_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[4] ),
    .A2(net494),
    .B1(net491),
    .B2(\digitop_pav2.pie_inst.fsm.pivot[5] ),
    .C1(_10986_),
    .X(_10987_));
 o221a_1 _15910_ (.A1(net1300),
    .A2(_09585_),
    .B1(net491),
    .B2(\digitop_pav2.pie_inst.fsm.pivot[5] ),
    .C1(_10987_),
    .X(_10988_));
 a2111o_1 _15911_ (.A1(net1300),
    .A2(_09585_),
    .B1(_10988_),
    .C1(\digitop_pav2.pie_inst.fsm.pivot[7] ),
    .D1(\digitop_pav2.pie_inst.fsm.pivot[8] ),
    .X(_10989_));
 nand2_2 _15912_ (.A(\digitop_pav2.pie_inst.fsm.past_ovf_b ),
    .B(_10989_),
    .Y(_10990_));
 and3_1 _15913_ (.A(\digitop_pav2.pie_inst.fsm.past_ovf_b ),
    .B(_10981_),
    .C(_10989_),
    .X(_10991_));
 and2_1 _15914_ (.A(_07145_),
    .B(\digitop_pav2.pie_inst.fsm.state[1] ),
    .X(_10992_));
 or2_1 _15915_ (.A(\digitop_pav2.pie_inst.fsm.pivot[4] ),
    .B(net495),
    .X(_10993_));
 o211a_1 _15916_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[1] ),
    .A2(_09576_),
    .B1(_10957_),
    .C1(\digitop_pav2.pie_inst.fsm.pivot[0] ),
    .X(_10994_));
 a221o_1 _15917_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[1] ),
    .A2(_09576_),
    .B1(_09583_),
    .B2(\digitop_pav2.pie_inst.fsm.pivot[2] ),
    .C1(_10994_),
    .X(_10995_));
 o221a_1 _15918_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[2] ),
    .A2(_09583_),
    .B1(_10949_),
    .B2(net1301),
    .C1(_10995_),
    .X(_10996_));
 a221o_1 _15919_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[4] ),
    .A2(net495),
    .B1(_10949_),
    .B2(net1301),
    .C1(_10996_),
    .X(_10997_));
 a22o_1 _15920_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[5] ),
    .A2(net493),
    .B1(_10993_),
    .B2(_10997_),
    .X(_10998_));
 o221a_1 _15921_ (.A1(net1300),
    .A2(net494),
    .B1(net493),
    .B2(\digitop_pav2.pie_inst.fsm.pivot[5] ),
    .C1(_10998_),
    .X(_10999_));
 a221o_1 _15922_ (.A1(net1300),
    .A2(net494),
    .B1(net491),
    .B2(\digitop_pav2.pie_inst.fsm.pivot[7] ),
    .C1(_10999_),
    .X(_11000_));
 o22a_1 _15923_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[8] ),
    .A2(_09585_),
    .B1(net491),
    .B2(\digitop_pav2.pie_inst.fsm.pivot[7] ),
    .X(_11001_));
 a22o_1 _15924_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[8] ),
    .A2(_09585_),
    .B1(_11000_),
    .B2(_11001_),
    .X(_11002_));
 nor2_1 _15925_ (.A(_07145_),
    .B(\digitop_pav2.pie_inst.fsm.state[1] ),
    .Y(_11003_));
 a21o_1 _15926_ (.A1(_11002_),
    .A2(_11003_),
    .B1(_10992_),
    .X(_11004_));
 and2_1 _15927_ (.A(_10991_),
    .B(_11004_),
    .X(\digitop_pav2.pie_inst.fsm.n_data_en ));
 a211o_1 _15928_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[12] ),
    .A2(net156),
    .B1(_08518_),
    .C1(_10507_),
    .X(\digitop_pav2.proc_ctrl_inst.cmdfsm.n_crc_eval ));
 or4_1 _15929_ (.A(net137),
    .B(net136),
    .C(net135),
    .D(net134),
    .X(_11005_));
 or3_1 _15930_ (.A(net130),
    .B(net133),
    .C(net119),
    .X(_11006_));
 or3_4 _15931_ (.A(net108),
    .B(_11005_),
    .C(_11006_),
    .X(net84));
 or4_1 _15932_ (.A(net111),
    .B(net112),
    .C(net113),
    .D(net114),
    .X(_11007_));
 or3_1 _15933_ (.A(net139),
    .B(net109),
    .C(net110),
    .X(_11008_));
 or3_4 _15934_ (.A(net138),
    .B(_11007_),
    .C(_11008_),
    .X(net85));
 a311o_1 _15935_ (.A1(_09393_),
    .A2(_09400_),
    .A3(_09403_),
    .B1(_09397_),
    .C1(_09389_),
    .X(_11009_));
 or4b_4 _15936_ (.A(net118),
    .B(net121),
    .C(net123),
    .D_N(_11009_),
    .X(net86));
 or4_1 _15937_ (.A(net128),
    .B(net129),
    .C(net131),
    .D(net132),
    .X(_11010_));
 a211o_1 _15938_ (.A1(_09403_),
    .A2(_09405_),
    .B1(_09389_),
    .C1(_09398_),
    .X(_11011_));
 or4b_4 _15939_ (.A(net124),
    .B(net125),
    .C(_11010_),
    .D_N(_11011_),
    .X(net87));
 a31o_1 _15940_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[7] ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_end_i ),
    .A3(_09592_),
    .B1(_09611_),
    .X(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.n_int_wr_bit ));
 o31a_1 _15941_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[7] ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[6] ),
    .A3(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[5] ),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_end_i ),
    .X(_11012_));
 a22o_1 _15942_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.form_end ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[0] ),
    .B1(_09592_),
    .B2(_11012_),
    .X(_11013_));
 or3_1 _15943_ (.A(_09603_),
    .B(_09611_),
    .C(_11013_),
    .X(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.n_int_wr_stb ));
 and4bb_1 _15944_ (.A_N(_09591_),
    .B_N(_09613_),
    .C(_09609_),
    .D(net1480),
    .X(_11014_));
 and2_1 _15945_ (.A(_09591_),
    .B(_11012_),
    .X(_11015_));
 and4_1 _15946_ (.A(net1480),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[2] ),
    .C(_09592_),
    .D(_09598_),
    .X(_11016_));
 or3_1 _15947_ (.A(_11014_),
    .B(_11015_),
    .C(_11016_),
    .X(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.n_int_rd_stb ));
 or2_1 _15948_ (.A(_09643_),
    .B(_09644_),
    .X(_11017_));
 or4b_1 _15949_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_int_wr_bit ),
    .B(_09645_),
    .C(_09646_),
    .D_N(_11017_),
    .X(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_int_wr_stb ));
 or4_1 _15950_ (.A(net188),
    .B(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[3] ),
    .C(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[2] ),
    .D(net531),
    .X(_11018_));
 o311a_1 _15951_ (.A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[1] ),
    .A2(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[0] ),
    .A3(_09557_),
    .B1(_11018_),
    .C1(_09552_),
    .X(_11019_));
 or3_1 _15952_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[1] ),
    .B(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[0] ),
    .C(_09554_),
    .X(_11020_));
 o211a_1 _15953_ (.A1(net188),
    .A2(_09540_),
    .B1(_09551_),
    .C1(_11020_),
    .X(_11021_));
 or3b_2 _15954_ (.A(_11019_),
    .B(_11021_),
    .C_N(_09548_),
    .X(_11022_));
 nor2_1 _15955_ (.A(net529),
    .B(_11022_),
    .Y(_11023_));
 inv_2 _15956_ (.A(_11023_),
    .Y(_11024_));
 or3b_1 _15957_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[2] ),
    .B(net190),
    .C_N(net191),
    .X(_11025_));
 or2_1 _15958_ (.A(_11023_),
    .B(_11025_),
    .X(_11026_));
 inv_2 _15959_ (.A(_11026_),
    .Y(_11027_));
 o211ai_1 _15960_ (.A1(_07123_),
    .A2(_09557_),
    .B1(_09560_),
    .C1(_09552_),
    .Y(_11028_));
 o21bai_1 _15961_ (.A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[1] ),
    .A2(_07123_),
    .B1_N(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[2] ),
    .Y(_11029_));
 a31o_1 _15962_ (.A1(net188),
    .A2(_07124_),
    .A3(_11029_),
    .B1(_09555_),
    .X(_11030_));
 o311a_1 _15963_ (.A1(net188),
    .A2(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[0] ),
    .A3(_10862_),
    .B1(_09554_),
    .C1(_09551_),
    .X(_11031_));
 o21ai_1 _15964_ (.A1(_07123_),
    .A2(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[2] ),
    .B1(_09556_),
    .Y(_11032_));
 a211o_1 _15965_ (.A1(_09552_),
    .A2(_11032_),
    .B1(_11031_),
    .C1(net529),
    .X(_11033_));
 a31oi_1 _15966_ (.A1(net529),
    .A2(_11028_),
    .A3(_11030_),
    .B1(_09547_),
    .Y(_11034_));
 and2b_1 _15967_ (.A_N(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[6] ),
    .B(_09547_),
    .X(_11035_));
 nor2_1 _15968_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[0] ),
    .B(_09543_),
    .Y(_11036_));
 nand2_1 _15969_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[2] ),
    .B(_09545_),
    .Y(_11037_));
 a211o_1 _15970_ (.A1(_11033_),
    .A2(_11034_),
    .B1(_11035_),
    .C1(_09545_),
    .X(_11038_));
 a31o_1 _15971_ (.A1(_09543_),
    .A2(_11037_),
    .A3(_11038_),
    .B1(_11036_),
    .X(_11039_));
 inv_2 _15972_ (.A(_11039_),
    .Y(_11040_));
 mux2_1 _15973_ (.A0(_08955_),
    .A1(_07043_),
    .S(\digitop_pav2.crc_inst.mctrl_data_end_ff ),
    .X(_11041_));
 mux2_2 _15974_ (.A0(_11040_),
    .A1(_11041_),
    .S(_09542_),
    .X(_11042_));
 nor2_1 _15975_ (.A(net531),
    .B(_11042_),
    .Y(_11043_));
 or2_1 _15976_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[1] ),
    .B(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[0] ),
    .X(_11044_));
 or2_2 _15977_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[2] ),
    .B(_11044_),
    .X(_11045_));
 inv_2 _15978_ (.A(_11045_),
    .Y(_11046_));
 a31o_1 _15979_ (.A1(_11022_),
    .A2(_11043_),
    .A3(_11046_),
    .B1(_11026_),
    .X(_11047_));
 nand2_1 _15980_ (.A(net529),
    .B(_11042_),
    .Y(_11048_));
 or4b_1 _15981_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[2] ),
    .B(_09537_),
    .C(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[1] ),
    .D_N(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[0] ),
    .X(_11049_));
 nand2_1 _15982_ (.A(net530),
    .B(_11049_),
    .Y(_11050_));
 xnor2_1 _15983_ (.A(_07125_),
    .B(_09546_),
    .Y(_11051_));
 a21oi_1 _15984_ (.A1(_07125_),
    .A2(_07126_),
    .B1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[0] ),
    .Y(_11052_));
 o211a_1 _15985_ (.A1(_07125_),
    .A2(_07126_),
    .B1(_09537_),
    .C1(_11052_),
    .X(_11053_));
 a21oi_1 _15986_ (.A1(_11051_),
    .A2(_11053_),
    .B1(_11050_),
    .Y(_11054_));
 nand2_1 _15987_ (.A(_11045_),
    .B(_11054_),
    .Y(_11055_));
 a21bo_1 _15988_ (.A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.n_data_valid ),
    .A2(_11046_),
    .B1_N(_11055_),
    .X(_11056_));
 and3b_1 _15989_ (.A_N(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[2] ),
    .B(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[0] ),
    .C(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[1] ),
    .X(_11057_));
 o211a_1 _15990_ (.A1(_11048_),
    .A2(_11056_),
    .B1(_11057_),
    .C1(_11024_),
    .X(_11058_));
 or4bb_1 _15991_ (.A(net189),
    .B(_11058_),
    .C_N(net191),
    .D_N(_11047_),
    .X(\digitop_pav2.fm0miller_inst.fm0x_ctrl.n_gand ));
 and3b_1 _15992_ (.A_N(net191),
    .B(net190),
    .C(net189),
    .X(_11059_));
 nand3b_1 _15993_ (.A_N(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[0] ),
    .B(net190),
    .C(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[2] ),
    .Y(_11060_));
 nand2_1 _15994_ (.A(net529),
    .B(_11045_),
    .Y(_11061_));
 nor2_1 _15995_ (.A(_11054_),
    .B(_11061_),
    .Y(_11062_));
 nor3b_2 _15996_ (.A(net191),
    .B(net190),
    .C_N(net189),
    .Y(_11063_));
 and3_1 _15997_ (.A(_11042_),
    .B(_11062_),
    .C(_11063_),
    .X(_11064_));
 a31o_1 _15998_ (.A1(_11043_),
    .A2(_11046_),
    .A3(_11059_),
    .B1(_11064_),
    .X(\digitop_pav2.fm0miller_inst.fm0x_ctrl.n_gor ));
 and2_1 _15999_ (.A(net159),
    .B(_07845_),
    .X(_11065_));
 a31o_1 _16000_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[1] ),
    .A2(_07056_),
    .A3(_07843_),
    .B1(_11065_),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_end ));
 nor3b_1 _16001_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[1] ),
    .B(net1310),
    .C_N(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[2] ),
    .Y(_11066_));
 a21oi_1 _16002_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[1] ),
    .A2(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[2] ),
    .B1(net1310),
    .Y(_11067_));
 a31o_1 _16003_ (.A1(net1826),
    .A2(_07848_),
    .A3(_11067_),
    .B1(_11065_),
    .X(_11068_));
 a21o_1 _16004_ (.A1(\digitop_pav2.access_inst.access_ctrl0.nvm_busy_i ),
    .A2(_07849_),
    .B1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_wr_stb ),
    .X(_11069_));
 or3_1 _16005_ (.A(net1310),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[2] ),
    .C(_07848_),
    .X(_11070_));
 inv_2 _16006_ (.A(_11070_),
    .Y(_11071_));
 a22o_1 _16007_ (.A1(net1310),
    .A2(_07844_),
    .B1(_11071_),
    .B2(net1826),
    .X(_11072_));
 or3_1 _16008_ (.A(_11068_),
    .B(_11069_),
    .C(_11072_),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_state[0] ));
 a21oi_1 _16009_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[0] ),
    .A2(net159),
    .B1(_07847_),
    .Y(_11073_));
 or4_1 _16010_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[1] ),
    .B(_07056_),
    .C(net1310),
    .D(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.ref_pulse_sync_o ),
    .X(_11074_));
 or4b_1 _16011_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[0] ),
    .B(net1310),
    .C(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[2] ),
    .D_N(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[1] ),
    .X(_11075_));
 o211a_1 _16012_ (.A1(_07056_),
    .A2(_07844_),
    .B1(_11074_),
    .C1(_11075_),
    .X(_11076_));
 or3b_1 _16013_ (.A(_11072_),
    .B(_11073_),
    .C_N(_11076_),
    .X(_11077_));
 nor2_1 _16014_ (.A(net1083),
    .B(_07898_),
    .Y(_11078_));
 xor2_1 _16015_ (.A(net1106),
    .B(\digitop_pav2.access_inst.access_check0.fg_i[8] ),
    .X(_11079_));
 xnor2_1 _16016_ (.A(net1114),
    .B(\digitop_pav2.cal_inst.calx_mux.dtest_trim_1_i ),
    .Y(_11080_));
 xor2_1 _16017_ (.A(net1110),
    .B(\digitop_pav2.cal_inst.calx_mux.dtest_trim_2_i ),
    .X(_11081_));
 xnor2_1 _16018_ (.A(net1098),
    .B(\digitop_pav2.access_inst.access_check0.fg_i[10] ),
    .Y(_11082_));
 o221ai_1 _16019_ (.A1(_07077_),
    .A2(net1323),
    .B1(\digitop_pav2.access_inst.access_check0.fg_i[13] ),
    .B2(_07083_),
    .C1(_11082_),
    .Y(_11083_));
 a221o_1 _16020_ (.A1(_07075_),
    .A2(\digitop_pav2.access_inst.access_check0.fg_i[1] ),
    .B1(\digitop_pav2.cal_inst.calx_mux.dtest_trim_0_i ),
    .B2(net1117),
    .C1(_11079_),
    .X(_11084_));
 a221o_1 _16021_ (.A1(net1123),
    .A2(_07096_),
    .B1(\digitop_pav2.access_inst.access_check0.fg_i[11] ),
    .B2(net1035),
    .C1(_11080_),
    .X(_11085_));
 a2bb2o_1 _16022_ (.A1_N(_07081_),
    .A2_N(\digitop_pav2.access_inst.access_check0.fg_i[11] ),
    .B1(\digitop_pav2.access_inst.access_check0.fg_i[9] ),
    .B2(_07080_),
    .X(_11086_));
 a221o_1 _16023_ (.A1(net1127),
    .A2(_07095_),
    .B1(net1323),
    .B2(_07077_),
    .C1(_11086_),
    .X(_11087_));
 or4_1 _16024_ (.A(_11083_),
    .B(_11084_),
    .C(_11085_),
    .D(_11087_),
    .X(_11088_));
 or4b_1 _16025_ (.A(_11078_),
    .B(_11081_),
    .C(_11088_),
    .D_N(_11065_),
    .X(_11089_));
 a22o_1 _16026_ (.A1(_07076_),
    .A2(\digitop_pav2.access_inst.access_check0.fg_i[3] ),
    .B1(_07117_),
    .B2(_07078_),
    .X(_11090_));
 a221o_1 _16027_ (.A1(_07083_),
    .A2(\digitop_pav2.access_inst.access_check0.fg_i[13] ),
    .B1(net1319),
    .B2(net1090),
    .C1(_11090_),
    .X(_11091_));
 nand2_1 _16028_ (.A(net1126),
    .B(\digitop_pav2.access_inst.access_check0.fg_i[2] ),
    .Y(_11092_));
 or2_1 _16029_ (.A(net1126),
    .B(\digitop_pav2.access_inst.access_check0.fg_i[2] ),
    .X(_11093_));
 nand2_1 _16030_ (.A(net1132),
    .B(net1324),
    .Y(_11094_));
 or2_1 _16031_ (.A(net1132),
    .B(net1324),
    .X(_11095_));
 a221o_1 _16032_ (.A1(_11092_),
    .A2(_11093_),
    .B1(_11094_),
    .B2(_11095_),
    .C1(_08104_),
    .X(_11096_));
 a211o_1 _16033_ (.A1(_07082_),
    .A2(net1318),
    .B1(_11091_),
    .C1(_11096_),
    .X(_11097_));
 a211o_1 _16034_ (.A1(net1083),
    .A2(_07898_),
    .B1(_11089_),
    .C1(_11097_),
    .X(_11098_));
 nand2b_1 _16035_ (.A_N(_11077_),
    .B(_11098_),
    .Y(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_state[1] ));
 a211o_1 _16036_ (.A1(_07115_),
    .A2(_11071_),
    .B1(_11073_),
    .C1(_11066_),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_state[2] ));
 or2_1 _16037_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[3] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_rd_stb ),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_state[3] ));
 mux2_1 _16038_ (.A0(\digitop_pav2.func_rr_erase ),
    .A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.rr_erase ),
    .S(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.tm_mbist_i ),
    .X(_11099_));
 and2_1 _16039_ (.A(net1494),
    .B(_11099_),
    .X(ff_erase));
 mux2_1 _16040_ (.A0(\digitop_pav2.func_rr_prog ),
    .A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.rr_prog ),
    .S(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.tm_mbist_i ),
    .X(_11100_));
 and2_1 _16041_ (.A(net1494),
    .B(_11100_),
    .X(ff_prog));
 nor2_1 _16042_ (.A(_00154_),
    .B(_00574_),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux_before_buf ));
 nand3_1 _16043_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk_before_buf ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.en_ctr ),
    .C(net514),
    .Y(_00155_));
 nand2b_1 _16044_ (.A_N(net1250),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div4_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_en.piex_clk_dis ));
 and2_1 _16045_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[1] ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[0] ),
    .X(_11101_));
 and3_1 _16046_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[3] ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[2] ),
    .C(_11101_),
    .X(_11102_));
 and2_1 _16047_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[4] ),
    .B(_11102_),
    .X(_11103_));
 and3_1 _16048_ (.A(net1827),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[4] ),
    .C(_11102_),
    .X(_11104_));
 inv_2 _16049_ (.A(net1828),
    .Y(_00161_));
 nand2_2 _16050_ (.A(_00237_),
    .B(\digitop_pav2.pie_inst.fsm.past_clk_i ),
    .Y(\digitop_pav2.pie_inst.en_ctr ));
 nand2_1 _16051_ (.A(_07843_),
    .B(_07848_),
    .Y(_11105_));
 and2_1 _16052_ (.A(net1310),
    .B(_11105_),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_end_stab_clk ));
 and2_1 _16053_ (.A(net1233),
    .B(\digitop_pav2.ack_inst.state_ff[0] ),
    .X(_00006_));
 and2b_1 _16054_ (.A_N(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.form_end ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[0] ),
    .X(_00012_));
 and2b_1 _16055_ (.A_N(net1481),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[0] ),
    .X(_00013_));
 and2_1 _16056_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[0] ),
    .B(_09626_),
    .X(_00011_));
 nor2_1 _16057_ (.A(_07121_),
    .B(_08504_),
    .Y(_00010_));
 and2_1 _16058_ (.A(\digitop_pav2.sec_inst.shift_out.st[2] ),
    .B(_08504_),
    .X(_00009_));
 nor2_1 _16059_ (.A(_07121_),
    .B(_08505_),
    .Y(_00008_));
 o22a_1 _16060_ (.A1(_09492_),
    .A2(_10761_),
    .B1(_10764_),
    .B2(_10760_),
    .X(_11106_));
 nor2_1 _16061_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.n_state[4] ),
    .B(_11106_),
    .Y(_11107_));
 or4_1 _16062_ (.A(\digitop_pav2.testctrl_pav2.inst_mode.tm_amux ),
    .B(_09463_),
    .C(_09482_),
    .D(_11107_),
    .X(_00162_));
 or4b_2 _16063_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[1] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[2] ),
    .C(_09633_),
    .D_N(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[0] ),
    .X(_11108_));
 and4b_1 _16064_ (.A_N(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[15] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[2] ),
    .C(_09635_),
    .D(_11108_),
    .X(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_prog ));
 and4_1 _16065_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[15] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[2] ),
    .C(_09635_),
    .D(_11108_),
    .X(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_erase ));
 o21a_1 _16066_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[5] ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[7] ),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_end_i ),
    .X(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_int_rd_stb ));
 or2_1 _16067_ (.A(\digitop_pav2.func_rnclk_en ),
    .B(\digitop_pav2.testctrl_pav2.inst_mode.tm_rnclkout ),
    .X(net80));
 a221o_1 _16068_ (.A1(net1483),
    .A2(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.nvm_calx_rd_stb_o ),
    .B1(_09166_),
    .B2(\digitop_pav2.sec_inst.ld_mem.st[0] ),
    .C1(_09167_),
    .X(_11109_));
 or4b_2 _16069_ (.A(\digitop_pav2.ack_inst.nvm_ack_rd_stb_o ),
    .B(_09162_),
    .C(_11109_),
    .D_N(_09163_),
    .X(\digitop_pav2.glue_inst.mbus_rd_en_o ));
 nor2_1 _16070_ (.A(_07839_),
    .B(net1778),
    .Y(_11110_));
 a211o_1 _16071_ (.A1(net1482),
    .A2(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.nvm_calx_wr_stb_o ),
    .B1(_09164_),
    .C1(_11110_),
    .X(\digitop_pav2.glue_inst.mbus_wr_en_o ));
 or3_1 _16072_ (.A(net1755),
    .B(_07058_),
    .C(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_replay_o ),
    .X(_11111_));
 o21ai_1 _16073_ (.A1(net1779),
    .A2(net1314),
    .B1(_08324_),
    .Y(\digitop_pav2.stadly_memctrl_wr_dt0_0.A ));
 and2_1 _16074_ (.A(net1482),
    .B(_11069_),
    .X(_11112_));
 nor2_1 _16075_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[1] ),
    .B(net1314),
    .Y(_11113_));
 a211o_1 _16076_ (.A1(net1324),
    .A2(net155),
    .B1(_11113_),
    .C1(_08293_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt1_0.A ));
 nor2_1 _16077_ (.A(net1804),
    .B(net1314),
    .Y(_11114_));
 a211o_1 _16078_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[1] ),
    .A2(net155),
    .B1(_11114_),
    .C1(_08259_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt2_0.A ));
 nor2_1 _16079_ (.A(net1801),
    .B(net1314),
    .Y(_11115_));
 a211o_1 _16080_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[2] ),
    .A2(net155),
    .B1(_11115_),
    .C1(_08153_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt3_0.A ));
 nor2_1 _16081_ (.A(net1799),
    .B(net1315),
    .Y(_11116_));
 a211o_1 _16082_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[3] ),
    .A2(net155),
    .B1(_11116_),
    .C1(_08171_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt4_0.A ));
 nor2_1 _16083_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[5] ),
    .B(net1315),
    .Y(_11117_));
 a211o_1 _16084_ (.A1(net1323),
    .A2(net155),
    .B1(_11117_),
    .C1(_08372_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt5_0.A ));
 nor2_1 _16085_ (.A(net1794),
    .B(net1315),
    .Y(_11118_));
 a311o_1 _16086_ (.A1(net1482),
    .A2(_07117_),
    .A3(_11069_),
    .B1(_11118_),
    .C1(_08225_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt6_0.A ));
 o21ai_1 _16087_ (.A1(net1784),
    .A2(net1314),
    .B1(_08341_),
    .Y(_11119_));
 a31o_1 _16088_ (.A1(net1482),
    .A2(_07116_),
    .A3(_11069_),
    .B1(net1785),
    .X(\digitop_pav2.stadly_memctrl_wr_dt7_0.A ));
 nor2_1 _16089_ (.A(net1787),
    .B(net1314),
    .Y(_11120_));
 a311o_1 _16090_ (.A1(net1482),
    .A2(\digitop_pav2.cal_inst.calx_mux.dtest_trim_2_i ),
    .A3(_11069_),
    .B1(_11120_),
    .C1(_08356_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt8_0.A ));
 nor2_1 _16091_ (.A(net1795),
    .B(net1314),
    .Y(_11121_));
 a211o_1 _16092_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[8] ),
    .A2(_11112_),
    .B1(_11121_),
    .C1(_08188_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt9_0.A ));
 nor2_1 _16093_ (.A(net1792),
    .B(net1314),
    .Y(_11122_));
 a211o_1 _16094_ (.A1(\digitop_pav2.access_inst.access_check0.fg_i[9] ),
    .A2(net155),
    .B1(_11122_),
    .C1(_08276_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt10_0.A ));
 nor2_1 _16095_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[11] ),
    .B(net1315),
    .Y(_11123_));
 a211o_1 _16096_ (.A1(net1797),
    .A2(net155),
    .B1(_11123_),
    .C1(_08387_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt11_0.A ));
 nor2_1 _16097_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[12] ),
    .B(net1315),
    .Y(_11124_));
 a211o_1 _16098_ (.A1(net1790),
    .A2(net155),
    .B1(_11124_),
    .C1(_08308_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt12_0.A ));
 nor2_1 _16099_ (.A(net1803),
    .B(net1314),
    .Y(_11125_));
 a211o_1 _16100_ (.A1(net1318),
    .A2(net155),
    .B1(_11125_),
    .C1(_08207_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt13_0.A ));
 nor2_1 _16101_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[14] ),
    .B(net1314),
    .Y(_11126_));
 a211o_1 _16102_ (.A1(net1788),
    .A2(_11112_),
    .B1(_11126_),
    .C1(_08399_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt14_0.A ));
 nor2_1 _16103_ (.A(net1786),
    .B(net1315),
    .Y(_11127_));
 a211o_1 _16104_ (.A1(_07899_),
    .A2(net155),
    .B1(_11127_),
    .C1(_08241_),
    .X(\digitop_pav2.stadly_memctrl_wr_dt15_0.A ));
 and2_2 _16105_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_mask ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_pre_clk_before_buf ));
 or2_1 _16106_ (.A(net500),
    .B(_09271_),
    .X(_11128_));
 a21oi_1 _16107_ (.A1(_09273_),
    .A2(_11128_),
    .B1(_00149_),
    .Y(_11129_));
 nand2_1 _16108_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[7].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Y(_11130_));
 xnor2_1 _16109_ (.A(_09250_),
    .B(_09273_),
    .Y(_11131_));
 mux2_1 _16110_ (.A0(_09883_),
    .A1(net515),
    .S(_09273_),
    .X(_11132_));
 xnor2_1 _16111_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .B(_09865_),
    .Y(_11133_));
 xnor2_1 _16112_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .B(net508),
    .Y(_11134_));
 xnor2_1 _16113_ (.A(_00146_),
    .B(net522),
    .Y(_11135_));
 or2_1 _16114_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[7].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .X(_11136_));
 a311o_1 _16115_ (.A1(_00149_),
    .A2(_09273_),
    .A3(_11128_),
    .B1(_11129_),
    .C1(_11133_),
    .X(_11137_));
 or3_1 _16116_ (.A(_11134_),
    .B(_11135_),
    .C(_11137_),
    .X(_11138_));
 xnor2_1 _16117_ (.A(_00151_),
    .B(_11132_),
    .Y(_11139_));
 xnor2_1 _16118_ (.A(_00150_),
    .B(_11131_),
    .Y(_11140_));
 mux2_1 _16119_ (.A0(_11130_),
    .A1(_11136_),
    .S(_09281_),
    .X(_11141_));
 or4_1 _16120_ (.A(_11138_),
    .B(_11139_),
    .C(_11140_),
    .D(_11141_),
    .X(_11142_));
 or3b_1 _16121_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk_before_buf ),
    .B(_09282_),
    .C_N(_11142_),
    .X(_11143_));
 nor2_1 _16122_ (.A(net508),
    .B(_10191_),
    .Y(_11144_));
 inv_2 _16123_ (.A(_11144_),
    .Y(_11145_));
 nand2_1 _16124_ (.A(net508),
    .B(_10191_),
    .Y(_11146_));
 mux2_1 _16125_ (.A0(_11145_),
    .A1(_11146_),
    .S(net511),
    .X(_11147_));
 mux2_1 _16126_ (.A0(net496),
    .A1(_09868_),
    .S(_11144_),
    .X(_11148_));
 nor2_1 _16127_ (.A(_11147_),
    .B(_11148_),
    .Y(_11149_));
 and3_1 _16128_ (.A(net505),
    .B(_09864_),
    .C(_11144_),
    .X(_11150_));
 a21oi_1 _16129_ (.A1(_09864_),
    .A2(_11144_),
    .B1(net505),
    .Y(_11151_));
 or2_1 _16130_ (.A(_11150_),
    .B(_11151_),
    .X(_11152_));
 nand2_2 _16131_ (.A(_11149_),
    .B(_11152_),
    .Y(_11153_));
 or2_1 _16132_ (.A(_11149_),
    .B(_11152_),
    .X(_11154_));
 and2_1 _16133_ (.A(_11153_),
    .B(_11154_),
    .X(_11155_));
 xnor2_1 _16134_ (.A(_00150_),
    .B(_11155_),
    .Y(_11156_));
 or3b_1 _16135_ (.A(net511),
    .B(_11144_),
    .C_N(_11146_),
    .X(_11157_));
 nand2_1 _16136_ (.A(_11147_),
    .B(_11157_),
    .Y(_11158_));
 nor2_1 _16137_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .B(_11158_),
    .Y(_11159_));
 xnor2_1 _16138_ (.A(net513),
    .B(_11135_),
    .Y(_11160_));
 xnor2_1 _16139_ (.A(_10191_),
    .B(_11134_),
    .Y(_11161_));
 or3_1 _16140_ (.A(_11159_),
    .B(_11160_),
    .C(_11161_),
    .X(_11162_));
 a211o_1 _16141_ (.A1(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .A2(_11158_),
    .B1(_11162_),
    .C1(_09282_),
    .X(_11163_));
 xnor2_1 _16142_ (.A(_00151_),
    .B(net519),
    .Y(_11164_));
 xnor2_1 _16143_ (.A(_11150_),
    .B(_11164_),
    .Y(_11165_));
 o21bai_1 _16144_ (.A1(_11153_),
    .A2(_11165_),
    .B1_N(_11163_),
    .Y(_11166_));
 or4_1 _16145_ (.A(net520),
    .B(net519),
    .C(_11150_),
    .D(_11153_),
    .X(_11167_));
 a221o_1 _16146_ (.A1(_11153_),
    .A2(_11165_),
    .B1(_11167_),
    .B2(_00153_),
    .C1(_11166_),
    .X(_11168_));
 a21oi_1 _16147_ (.A1(net496),
    .A2(_11147_),
    .B1(_11149_),
    .Y(_11169_));
 xnor2_1 _16148_ (.A(_00149_),
    .B(_11169_),
    .Y(_11170_));
 a21boi_1 _16149_ (.A1(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .A2(_11167_),
    .B1_N(_11136_),
    .Y(_11171_));
 or4_1 _16150_ (.A(_11156_),
    .B(_11168_),
    .C(_11170_),
    .D(_11171_),
    .X(_11172_));
 nor2_1 _16151_ (.A(_10192_),
    .B(_11147_),
    .Y(_11173_));
 xnor2_1 _16152_ (.A(_11148_),
    .B(_11173_),
    .Y(_11174_));
 xnor2_1 _16153_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .B(_11174_),
    .Y(_11175_));
 o211a_1 _16154_ (.A1(net514),
    .A2(_09921_),
    .B1(_11145_),
    .C1(net501),
    .X(_11176_));
 o311a_1 _16155_ (.A1(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .A2(_11173_),
    .A3(_11176_),
    .B1(_11134_),
    .C1(_11160_),
    .X(_11177_));
 a21o_1 _16156_ (.A1(_10193_),
    .A2(_11149_),
    .B1(_11152_),
    .X(_11178_));
 o21a_1 _16157_ (.A1(_10192_),
    .A2(_11153_),
    .B1(_11178_),
    .X(_11179_));
 xnor2_1 _16158_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .B(_11179_),
    .Y(_11180_));
 and4_1 _16159_ (.A(_09282_),
    .B(_11175_),
    .C(_11177_),
    .D(_11180_),
    .X(_11181_));
 or3_1 _16160_ (.A(_10192_),
    .B(_11153_),
    .C(_11165_),
    .X(_11182_));
 o21ai_1 _16161_ (.A1(_10192_),
    .A2(_11153_),
    .B1(_11165_),
    .Y(_11183_));
 o21ai_1 _16162_ (.A1(_10192_),
    .A2(_11167_),
    .B1(_11130_),
    .Y(_11184_));
 and4_1 _16163_ (.A(_11181_),
    .B(_11182_),
    .C(_11183_),
    .D(_11184_),
    .X(_11185_));
 nand3b_1 _16164_ (.A_N(_11185_),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk_before_buf ),
    .C(_11172_),
    .Y(_11186_));
 a21o_1 _16165_ (.A1(_11143_),
    .A2(_11186_),
    .B1(_00154_),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_gen_cg.enable ));
 and3_2 _16166_ (.A(\digitop_pav2.cal_inst.calx_clk_o ),
    .B(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .C(\digitop_pav2.clkx_cp_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_merge.merge_clk ));
 and2_2 _16167_ (.A(\digitop_pav2.clkx_cp_clk ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.rngx_pup_clk_i ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_sel.rngx_clk ));
 o21a_1 _16168_ (.A1(\digitop_pav2.testctrl_pav2.inst_mode.tm_anafunc ),
    .A2(net1),
    .B1(_07113_),
    .X(_11187_));
 a211o_2 _16169_ (.A1(net1503),
    .A2(\digitop_pav2.testctrl_pav2.inst_mode.tm_digfunc ),
    .B1(_11187_),
    .C1(net1483),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_i ));
 xor2_1 _16170_ (.A(\digitop_pav2.rng_inst.rng_trngx_pav2.neg_data ),
    .B(\digitop_pav2.rng_inst.rng_trngx_pav2.pos_data ),
    .X(\digitop_pav2.rng_inst.rng_trngx_pav2.xor_data ));
 a21oi_1 _16171_ (.A1(net1290),
    .A2(net1188),
    .B1(net1295),
    .Y(_11188_));
 o21ai_1 _16172_ (.A1(_07294_),
    .A2(_11188_),
    .B1(_10465_),
    .Y(\digitop_pav2.proc_ctrl_inst.cmdfsm.cg_en_out2 ));
 or2_1 _16173_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_cgen.en_g_sec_i ),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_cgen.fg_tc_rx_i ),
    .X(_11189_));
 a221o_1 _16174_ (.A1(_07153_),
    .A2(_09024_),
    .B1(_11189_),
    .B2(net1294),
    .C1(_10490_),
    .X(\digitop_pav2.proc_ctrl_inst.cmdfsm.cg_en_out1 ));
 and2b_1 _16175_ (.A_N(net1807),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmd_abort_b ),
    .X(\digitop_pav2.proc_ctrl_inst.cmd.rst_b_i ));
 and2_2 _16176_ (.A(\digitop_pav2.pie_inst.en_ctr_fix ),
    .B(net1225),
    .X(\digitop_pav2.pie_inst.ctr.en_ctr_i ));
 and2_1 _16177_ (.A(_07061_),
    .B(_10318_),
    .X(\digitop_pav2.memctrl_inst.n_prog ));
 and2_1 _16178_ (.A(net1083),
    .B(_10318_),
    .X(\digitop_pav2.memctrl_inst.n_erase ));
 nor2_1 _16179_ (.A(_07047_),
    .B(net1398),
    .Y(\digitop_pav2.invent_inst.s2_s_o ));
 and2_1 _16180_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_r_ff_i ),
    .B(net1453),
    .X(\digitop_pav2.invent_inst.s2_r_o ));
 nor2_1 _16181_ (.A(_07046_),
    .B(net1398),
    .Y(\digitop_pav2.invent_inst.s3_s_o ));
 and2_1 _16182_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_r_ff_i ),
    .B(net1453),
    .X(\digitop_pav2.invent_inst.s3_r_o ));
 and2_1 _16183_ (.A(\digitop_pav2.invent_inst.sl_s_ff ),
    .B(net1452),
    .X(\digitop_pav2.invent_inst.sl_s_o ));
 and2_1 _16184_ (.A(\digitop_pav2.invent_inst.sl_r_ff ),
    .B(net1451),
    .X(\digitop_pav2.invent_inst.sl_r_o ));
 and3_2 _16185_ (.A(net1503),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.ref_pulse_sync_o ),
    .C(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.rp_ff[0] ),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk_dftmux.dft_rp_and ));
 or2_1 _16186_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.end_stab_clk_i ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.stab_clk_dis ),
    .X(_00133_));
 and2_2 _16187_ (.A(net1482),
    .B(clk_i),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.aux_clk ));
 and2_1 _16188_ (.A(\digitop_pav2.boot_inst.boot_ctrl0.state[0] ),
    .B(net1400),
    .X(_00007_));
 mux2_1 _16189_ (.A0(\digitop_pav2.func_rr_read ),
    .A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.rr_read ),
    .S(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.tm_mbist_i ),
    .X(_11190_));
 and2_1 _16190_ (.A(net68),
    .B(_11190_),
    .X(net107));
 and2_1 _16191_ (.A(net68),
    .B(_11099_),
    .X(net104));
 and2_1 _16192_ (.A(net68),
    .B(_11100_),
    .X(net106));
 or4_1 _16193_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[2] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[3] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[1] ),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.reg_wr_en ),
    .X(_00353_));
 o21ba_1 _16194_ (.A1(sl_set_ff2),
    .A2(\digitop_pav2.sl_i ),
    .B1_N(net1835),
    .X(_00354_));
 o21ba_1 _16195_ (.A1(s3_set_ff2),
    .A2(\digitop_pav2.s3_i ),
    .B1_N(net1830),
    .X(_00355_));
 o21ba_1 _16196_ (.A1(s2_set_ff2),
    .A2(\digitop_pav2.s2_i ),
    .B1_N(net1833),
    .X(_00356_));
 and2_1 _16197_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[4] ),
    .B(_10743_),
    .X(_11191_));
 nand2_1 _16198_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[4] ),
    .B(_10743_),
    .Y(_11192_));
 nor2_2 _16199_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[4] ),
    .B(net398),
    .Y(_11193_));
 nor2_4 _16200_ (.A(_11191_),
    .B(_11193_),
    .Y(_11194_));
 nor2_1 _16201_ (.A(net185),
    .B(_07110_),
    .Y(_11195_));
 nand2_1 _16202_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_9.Y ),
    .B(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_9.Y ),
    .Y(_11196_));
 a21oi_4 _16203_ (.A1(net417),
    .A2(_11196_),
    .B1(_11194_),
    .Y(_11197_));
 nand2_2 _16204_ (.A(net468),
    .B(_11196_),
    .Y(_11198_));
 nand2_1 _16205_ (.A(_07105_),
    .B(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[0] ),
    .Y(_11199_));
 nor2_1 _16206_ (.A(_07106_),
    .B(_11199_),
    .Y(_11200_));
 nor2_1 _16207_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[0] ),
    .Y(_11201_));
 nand2_1 _16208_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[2] ),
    .B(net404),
    .Y(_11202_));
 o2bb2a_1 _16209_ (.A1_N(_11191_),
    .A2_N(_11202_),
    .B1(net364),
    .B2(_07516_),
    .X(_11203_));
 and3_1 _16210_ (.A(_11197_),
    .B(_11198_),
    .C(_11203_),
    .X(_11204_));
 nor2_1 _16211_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[2] ),
    .B(_11199_),
    .Y(_11205_));
 or2_1 _16212_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[2] ),
    .B(_11199_),
    .X(_11206_));
 and2_2 _16213_ (.A(_07106_),
    .B(net404),
    .X(_11207_));
 nand2_1 _16214_ (.A(_07106_),
    .B(_11201_),
    .Y(_11208_));
 a22o_1 _16215_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[13] ),
    .A2(net362),
    .B1(net395),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[13] ),
    .X(_11209_));
 nand2_2 _16216_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[0] ),
    .Y(_11210_));
 nor2_1 _16217_ (.A(_07106_),
    .B(_11210_),
    .Y(_11211_));
 or2_2 _16218_ (.A(_07105_),
    .B(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[0] ),
    .X(_11212_));
 nor2_1 _16219_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[2] ),
    .B(_11212_),
    .Y(_11213_));
 or2_1 _16220_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[2] ),
    .B(_11212_),
    .X(_11214_));
 nor2_1 _16221_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[2] ),
    .B(_11210_),
    .Y(_11215_));
 or2_1 _16222_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[2] ),
    .B(_11210_),
    .X(_11216_));
 nor2_1 _16223_ (.A(_07106_),
    .B(_11212_),
    .Y(_11217_));
 a221o_1 _16224_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[5] ),
    .A2(net404),
    .B1(net389),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[5] ),
    .C1(net396),
    .X(_11218_));
 a22o_1 _16225_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[5] ),
    .A2(net361),
    .B1(net355),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[5] ),
    .X(_11219_));
 a221o_1 _16226_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[5] ),
    .A2(net365),
    .B1(net390),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[5] ),
    .C1(_11219_),
    .X(_11220_));
 a211o_1 _16227_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[5] ),
    .A2(net357),
    .B1(_11218_),
    .C1(_11220_),
    .X(_11221_));
 or2_1 _16228_ (.A(net439),
    .B(net426),
    .X(_11222_));
 or3_4 _16229_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[0] ),
    .B(_07521_),
    .C(net402),
    .X(_11223_));
 nor2_1 _16230_ (.A(net469),
    .B(_11223_),
    .Y(_11224_));
 or2_1 _16231_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[5] ),
    .B(net392),
    .X(_11225_));
 a32oi_1 _16232_ (.A1(_11221_),
    .A2(net351),
    .A3(_11225_),
    .B1(_11209_),
    .B2(net445),
    .Y(_11226_));
 a32o_1 _16233_ (.A1(_11221_),
    .A2(net351),
    .A3(_11225_),
    .B1(_11209_),
    .B2(net444),
    .X(_11227_));
 a22o_2 _16234_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[11] ),
    .A2(net360),
    .B1(net395),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[11] ),
    .X(_11228_));
 a221o_1 _16235_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[3] ),
    .A2(net365),
    .B1(net403),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[3] ),
    .C1(net396),
    .X(_11229_));
 a22o_1 _16236_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[3] ),
    .A2(net390),
    .B1(net356),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[3] ),
    .X(_11230_));
 a221o_1 _16237_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[3] ),
    .A2(net361),
    .B1(net388),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[3] ),
    .C1(_11230_),
    .X(_11231_));
 a211o_1 _16238_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[3] ),
    .A2(net354),
    .B1(_11229_),
    .C1(_11231_),
    .X(_11232_));
 or2_1 _16239_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[3] ),
    .B(net392),
    .X(_11233_));
 a32oi_1 _16240_ (.A1(net350),
    .A2(_11232_),
    .A3(_11233_),
    .B1(_11228_),
    .B2(net444),
    .Y(_11234_));
 a32o_1 _16241_ (.A1(net350),
    .A2(_11232_),
    .A3(_11233_),
    .B1(_11228_),
    .B2(net450),
    .X(_11235_));
 a22o_1 _16242_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[9] ),
    .A2(net363),
    .B1(net397),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[9] ),
    .X(_11236_));
 a22o_1 _16243_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[1] ),
    .A2(net361),
    .B1(net356),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[1] ),
    .X(_11237_));
 a221o_1 _16244_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[1] ),
    .A2(net403),
    .B1(net388),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[1] ),
    .C1(net396),
    .X(_11238_));
 a221o_1 _16245_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[1] ),
    .A2(net365),
    .B1(net390),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[1] ),
    .C1(_11238_),
    .X(_11239_));
 a211o_2 _16246_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[1] ),
    .A2(net354),
    .B1(_11237_),
    .C1(_11239_),
    .X(_11240_));
 or2_1 _16247_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[1] ),
    .B(net393),
    .X(_11241_));
 a32oi_4 _16248_ (.A1(net350),
    .A2(_11240_),
    .A3(_11241_),
    .B1(_11236_),
    .B2(net444),
    .Y(_11242_));
 a32o_1 _16249_ (.A1(net350),
    .A2(_11240_),
    .A3(_11241_),
    .B1(_11236_),
    .B2(net444),
    .X(_11243_));
 a22o_1 _16250_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[8] ),
    .A2(net360),
    .B1(net395),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[8] ),
    .X(_11244_));
 o21a_1 _16251_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[0] ),
    .A2(_07106_),
    .B1(net403),
    .X(_11245_));
 a221o_1 _16252_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[0] ),
    .A2(net390),
    .B1(net388),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ),
    .C1(_11245_),
    .X(_11246_));
 a22o_1 _16253_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[0] ),
    .A2(net365),
    .B1(net361),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[0] ),
    .X(_11247_));
 a221o_1 _16254_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[0] ),
    .A2(net356),
    .B1(net355),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[0] ),
    .C1(_11247_),
    .X(_11248_));
 o221a_1 _16255_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[0] ),
    .A2(net394),
    .B1(_11246_),
    .B2(_11248_),
    .C1(net353),
    .X(_11249_));
 a21oi_1 _16256_ (.A1(net449),
    .A2(_11244_),
    .B1(_11249_),
    .Y(_11250_));
 and2_1 _16257_ (.A(_11243_),
    .B(net236),
    .X(_11251_));
 nand2_4 _16258_ (.A(net288),
    .B(net235),
    .Y(_11252_));
 a22o_1 _16259_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[10] ),
    .A2(net360),
    .B1(net395),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[10] ),
    .X(_11253_));
 a221o_1 _16260_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[2] ),
    .A2(net364),
    .B1(net403),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[2] ),
    .C1(net396),
    .X(_11254_));
 a22o_1 _16261_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ),
    .A2(net390),
    .B1(net388),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[2] ),
    .X(_11255_));
 a221o_1 _16262_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[2] ),
    .A2(net361),
    .B1(net356),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[2] ),
    .C1(_11255_),
    .X(_11256_));
 a211o_1 _16263_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[2] ),
    .A2(net354),
    .B1(_11254_),
    .C1(_11256_),
    .X(_11257_));
 or2_1 _16264_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[2] ),
    .B(net392),
    .X(_11258_));
 a32o_2 _16265_ (.A1(net353),
    .A2(_11257_),
    .A3(_11258_),
    .B1(_11253_),
    .B2(net449),
    .X(_11259_));
 clkinv_4 _16266_ (.A(net287),
    .Y(_11260_));
 nor2_4 _16267_ (.A(net235),
    .B(net287),
    .Y(_11261_));
 or2_4 _16268_ (.A(net235),
    .B(net287),
    .X(_11262_));
 a21oi_2 _16269_ (.A1(_11252_),
    .A2(_11262_),
    .B1(net246),
    .Y(_11263_));
 or2_4 _16270_ (.A(net238),
    .B(net235),
    .X(_11264_));
 nand2_1 _16271_ (.A(net244),
    .B(_11252_),
    .Y(_11265_));
 nor2_1 _16272_ (.A(_11261_),
    .B(_11265_),
    .Y(_11266_));
 a22o_1 _16273_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[12] ),
    .A2(net362),
    .B1(_11207_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[12] ),
    .X(_11267_));
 a22o_1 _16274_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[4] ),
    .A2(net365),
    .B1(net355),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[4] ),
    .X(_11268_));
 a221o_1 _16275_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[4] ),
    .A2(net404),
    .B1(net357),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[4] ),
    .C1(net396),
    .X(_11269_));
 a221o_1 _16276_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[4] ),
    .A2(net361),
    .B1(net390),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[4] ),
    .C1(_11269_),
    .X(_11270_));
 a211o_1 _16277_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[4] ),
    .A2(net389),
    .B1(_11268_),
    .C1(_11270_),
    .X(_11271_));
 or2_1 _16278_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[4] ),
    .B(net392),
    .X(_11272_));
 a32oi_1 _16279_ (.A1(net350),
    .A2(_11271_),
    .A3(_11272_),
    .B1(_11267_),
    .B2(net444),
    .Y(_11273_));
 a32o_1 _16280_ (.A1(net350),
    .A2(_11271_),
    .A3(_11272_),
    .B1(_11267_),
    .B2(net445),
    .X(_11274_));
 nor2_2 _16281_ (.A(net288),
    .B(net235),
    .Y(_11275_));
 nor2_2 _16282_ (.A(net235),
    .B(_11260_),
    .Y(_11276_));
 or2_4 _16283_ (.A(net236),
    .B(_11260_),
    .X(_11277_));
 nand2_2 _16284_ (.A(net289),
    .B(_11276_),
    .Y(_11278_));
 nand2_1 _16285_ (.A(net236),
    .B(_11260_),
    .Y(_11279_));
 nor2_2 _16286_ (.A(net289),
    .B(net287),
    .Y(_11280_));
 nand2_4 _16287_ (.A(net288),
    .B(_11260_),
    .Y(_11281_));
 nand2_4 _16288_ (.A(net200),
    .B(_11281_),
    .Y(_11282_));
 nor2_1 _16289_ (.A(_11251_),
    .B(_11275_),
    .Y(_11283_));
 or2_2 _16290_ (.A(_11251_),
    .B(_11275_),
    .X(_11284_));
 nor2_1 _16291_ (.A(net287),
    .B(_11284_),
    .Y(_11285_));
 nand2_1 _16292_ (.A(_11252_),
    .B(_11282_),
    .Y(_11286_));
 and2_2 _16293_ (.A(net235),
    .B(net287),
    .X(_11287_));
 nand2_4 _16294_ (.A(net236),
    .B(net287),
    .Y(_11288_));
 nor2_2 _16295_ (.A(_11243_),
    .B(_11259_),
    .Y(_11289_));
 nand2_4 _16296_ (.A(net289),
    .B(_11260_),
    .Y(_11290_));
 nor2_1 _16297_ (.A(net288),
    .B(_11262_),
    .Y(_11291_));
 nand2_2 _16298_ (.A(net289),
    .B(_11261_),
    .Y(_11292_));
 nor2_2 _16299_ (.A(net289),
    .B(_11260_),
    .Y(_11293_));
 nand2_2 _16300_ (.A(net288),
    .B(net287),
    .Y(_11294_));
 nand2_1 _16301_ (.A(_11252_),
    .B(_11294_),
    .Y(_11295_));
 nand2_2 _16302_ (.A(_11260_),
    .B(_11284_),
    .Y(_11296_));
 nand2_1 _16303_ (.A(_11278_),
    .B(_11286_),
    .Y(_11297_));
 o21a_1 _16304_ (.A1(net240),
    .A2(_11297_),
    .B1(net233),
    .X(_11298_));
 a22o_1 _16305_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[14] ),
    .A2(net363),
    .B1(net397),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[14] ),
    .X(_11299_));
 a22o_1 _16306_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[6] ),
    .A2(net356),
    .B1(net388),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[6] ),
    .X(_11300_));
 a221o_1 _16307_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[6] ),
    .A2(net403),
    .B1(net390),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[6] ),
    .C1(net396),
    .X(_11301_));
 a221o_1 _16308_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[6] ),
    .A2(net365),
    .B1(net361),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[6] ),
    .C1(_11301_),
    .X(_11302_));
 a211o_1 _16309_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[6] ),
    .A2(net354),
    .B1(_11300_),
    .C1(_11302_),
    .X(_11303_));
 or2_1 _16310_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[6] ),
    .B(net393),
    .X(_11304_));
 a32oi_1 _16311_ (.A1(net351),
    .A2(_11303_),
    .A3(_11304_),
    .B1(_11299_),
    .B2(net445),
    .Y(_11305_));
 a32o_1 _16312_ (.A1(net351),
    .A2(_11303_),
    .A3(_11304_),
    .B1(_11299_),
    .B2(net444),
    .X(_11306_));
 nor2_1 _16313_ (.A(net238),
    .B(_11290_),
    .Y(_11307_));
 nand2_2 _16314_ (.A(_11252_),
    .B(net287),
    .Y(_11308_));
 inv_2 _16315_ (.A(_11308_),
    .Y(_11309_));
 or2_2 _16316_ (.A(_11275_),
    .B(_11308_),
    .X(_11310_));
 nor2_1 _16317_ (.A(net245),
    .B(_11289_),
    .Y(_11311_));
 nand2_2 _16318_ (.A(net238),
    .B(_11290_),
    .Y(_11312_));
 nor2_1 _16319_ (.A(_11242_),
    .B(_11288_),
    .Y(_11313_));
 nand2_1 _16320_ (.A(net288),
    .B(_11287_),
    .Y(_11314_));
 nand2_1 _16321_ (.A(net200),
    .B(_11310_),
    .Y(_11315_));
 or2_1 _16322_ (.A(_11312_),
    .B(_11315_),
    .X(_11316_));
 nand2_1 _16323_ (.A(_11264_),
    .B(net222),
    .Y(_11317_));
 nor2_1 _16324_ (.A(_11307_),
    .B(_11317_),
    .Y(_11318_));
 nor2_1 _16325_ (.A(net246),
    .B(_11308_),
    .Y(_11319_));
 nor2_2 _16326_ (.A(net246),
    .B(net288),
    .Y(_11320_));
 nand2_1 _16327_ (.A(net237),
    .B(net289),
    .Y(_11321_));
 o22a_1 _16328_ (.A1(net244),
    .A2(_11308_),
    .B1(_11320_),
    .B2(net200),
    .X(_11322_));
 o2bb2a_1 _16329_ (.A1_N(_11316_),
    .A2_N(_11318_),
    .B1(_11322_),
    .B2(net222),
    .X(_11323_));
 o21a_1 _16330_ (.A1(_11263_),
    .A2(_11266_),
    .B1(_11298_),
    .X(_11324_));
 a211o_1 _16331_ (.A1(net231),
    .A2(_11297_),
    .B1(_11263_),
    .C1(_11266_),
    .X(_11325_));
 nand2_1 _16332_ (.A(net285),
    .B(_11325_),
    .Y(_11326_));
 o22a_1 _16333_ (.A1(net285),
    .A2(_11323_),
    .B1(_11324_),
    .B2(_11326_),
    .X(_11327_));
 nand2_1 _16334_ (.A(net247),
    .B(net288),
    .Y(_11328_));
 nand2_4 _16335_ (.A(net245),
    .B(_11288_),
    .Y(_11329_));
 inv_2 _16336_ (.A(_11329_),
    .Y(_11330_));
 nand2_2 _16337_ (.A(net289),
    .B(_11287_),
    .Y(_11331_));
 nand2_1 _16338_ (.A(_11328_),
    .B(_11329_),
    .Y(_11332_));
 a221o_1 _16339_ (.A1(_11235_),
    .A2(_11275_),
    .B1(_11292_),
    .B2(_11332_),
    .C1(_11263_),
    .X(_11333_));
 nand2_1 _16340_ (.A(_11252_),
    .B(_11281_),
    .Y(_11334_));
 nand2_1 _16341_ (.A(net245),
    .B(_11278_),
    .Y(_11335_));
 o221a_1 _16342_ (.A1(net245),
    .A2(_11285_),
    .B1(_11334_),
    .B2(_11335_),
    .C1(net225),
    .X(_11336_));
 a211o_1 _16343_ (.A1(net231),
    .A2(_11333_),
    .B1(_11336_),
    .C1(net283),
    .X(_11337_));
 nor2_1 _16344_ (.A(net289),
    .B(net235),
    .Y(_11338_));
 or2_2 _16345_ (.A(net289),
    .B(net236),
    .X(_11339_));
 nor2_2 _16346_ (.A(_11260_),
    .B(_11338_),
    .Y(_11340_));
 or2_1 _16347_ (.A(net244),
    .B(_11340_),
    .X(_11341_));
 nand2_1 _16348_ (.A(net238),
    .B(net235),
    .Y(_11342_));
 nand2_1 _16349_ (.A(net238),
    .B(_11262_),
    .Y(_11343_));
 o21ai_2 _16350_ (.A1(_11340_),
    .A2(_11343_),
    .B1(net229),
    .Y(_11344_));
 inv_2 _16351_ (.A(_11344_),
    .Y(_11345_));
 nand2_1 _16352_ (.A(net242),
    .B(_11276_),
    .Y(_11346_));
 nor2_1 _16353_ (.A(_11289_),
    .B(_11293_),
    .Y(_11347_));
 nand2_1 _16354_ (.A(_11290_),
    .B(_11294_),
    .Y(_11348_));
 o211a_1 _16355_ (.A1(_11261_),
    .A2(_11348_),
    .B1(_11342_),
    .C1(net222),
    .X(_11349_));
 a311o_1 _16356_ (.A1(_11328_),
    .A2(_11345_),
    .A3(_11346_),
    .B1(_11349_),
    .C1(net284),
    .X(_11350_));
 a22o_1 _16357_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[15] ),
    .A2(net363),
    .B1(net397),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[15] ),
    .X(_11351_));
 a22o_1 _16358_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[7] ),
    .A2(net360),
    .B1(net354),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ),
    .X(_11352_));
 a221o_1 _16359_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[7] ),
    .A2(net403),
    .B1(net391),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ),
    .C1(net395),
    .X(_11353_));
 a221o_1 _16360_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[7] ),
    .A2(net364),
    .B1(net388),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ),
    .C1(_11353_),
    .X(_11354_));
 a211o_1 _16361_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ),
    .A2(net356),
    .B1(_11352_),
    .C1(_11354_),
    .X(_11355_));
 or2_1 _16362_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[7] ),
    .B(net393),
    .X(_11356_));
 a32oi_4 _16363_ (.A1(net350),
    .A2(_11355_),
    .A3(_11356_),
    .B1(_11351_),
    .B2(net446),
    .Y(_11357_));
 a32o_1 _16364_ (.A1(net350),
    .A2(_11355_),
    .A3(_11356_),
    .B1(_11351_),
    .B2(net444),
    .X(_11358_));
 a31o_1 _16365_ (.A1(net252),
    .A2(_11337_),
    .A3(_11350_),
    .B1(net281),
    .X(_11359_));
 a21oi_1 _16366_ (.A1(net249),
    .A2(_11327_),
    .B1(_11359_),
    .Y(_11360_));
 a31o_4 _16367_ (.A1(net462),
    .A2(_07105_),
    .A3(_07106_),
    .B1(net353),
    .X(_11361_));
 inv_2 _16368_ (.A(_11361_),
    .Y(_11362_));
 nand2_1 _16369_ (.A(_11252_),
    .B(_11277_),
    .Y(_11363_));
 nand2_1 _16370_ (.A(net236),
    .B(_11280_),
    .Y(_11364_));
 and3_1 _16371_ (.A(net243),
    .B(_11278_),
    .C(_11364_),
    .X(_11365_));
 nor2_1 _16372_ (.A(net244),
    .B(_11310_),
    .Y(_11366_));
 nand2_1 _16373_ (.A(net242),
    .B(net287),
    .Y(_11367_));
 nand2_1 _16374_ (.A(net247),
    .B(_11281_),
    .Y(_11368_));
 nor2_1 _16375_ (.A(net241),
    .B(_11280_),
    .Y(_11369_));
 nand2_1 _16376_ (.A(_11264_),
    .B(_11368_),
    .Y(_11370_));
 o32a_1 _16377_ (.A1(net230),
    .A2(_11365_),
    .A3(_11366_),
    .B1(_11370_),
    .B2(_11344_),
    .X(_11371_));
 nor2_1 _16378_ (.A(_11293_),
    .B(_11342_),
    .Y(_11372_));
 and3_1 _16379_ (.A(net244),
    .B(net200),
    .C(_11308_),
    .X(_11373_));
 o21a_1 _16380_ (.A1(_11372_),
    .A2(_11373_),
    .B1(net230),
    .X(_11374_));
 or2_1 _16381_ (.A(net239),
    .B(_11296_),
    .X(_11375_));
 nand2_1 _16382_ (.A(net239),
    .B(_11293_),
    .Y(_11376_));
 a31o_1 _16383_ (.A1(net223),
    .A2(_11375_),
    .A3(_11376_),
    .B1(net282),
    .X(_11377_));
 o22a_1 _16384_ (.A1(net284),
    .A2(_11371_),
    .B1(_11374_),
    .B2(_11377_),
    .X(_11378_));
 nor2_2 _16385_ (.A(net240),
    .B(_11293_),
    .Y(_11379_));
 nand2_1 _16386_ (.A(net242),
    .B(_11294_),
    .Y(_11380_));
 and2_1 _16387_ (.A(_11296_),
    .B(_11379_),
    .X(_11381_));
 and3_1 _16388_ (.A(net240),
    .B(_11288_),
    .C(_11292_),
    .X(_11382_));
 o21ai_1 _16389_ (.A1(_11381_),
    .A2(_11382_),
    .B1(net232),
    .Y(_11383_));
 and3_1 _16390_ (.A(_11262_),
    .B(_11281_),
    .C(_11332_),
    .X(_11384_));
 o311a_1 _16391_ (.A1(net232),
    .A2(_11319_),
    .A3(_11384_),
    .B1(_11383_),
    .C1(net283),
    .X(_11385_));
 or2_1 _16392_ (.A(_11251_),
    .B(_11282_),
    .X(_11386_));
 a21o_1 _16393_ (.A1(net240),
    .A2(_11386_),
    .B1(net225),
    .X(_11387_));
 or2_1 _16394_ (.A(_11332_),
    .B(_11387_),
    .X(_11388_));
 a2111o_1 _16395_ (.A1(net241),
    .A2(_11331_),
    .B1(_11313_),
    .C1(_11291_),
    .D1(net231),
    .X(_11389_));
 a31o_1 _16396_ (.A1(net285),
    .A2(_11388_),
    .A3(_11389_),
    .B1(net252),
    .X(_11390_));
 o221a_1 _16397_ (.A1(net249),
    .A2(_11378_),
    .B1(_11385_),
    .B2(_11390_),
    .C1(net281),
    .X(_11391_));
 or3_4 _16398_ (.A(_11360_),
    .B(_11362_),
    .C(_11391_),
    .X(_11392_));
 nor2_2 _16399_ (.A(_07092_),
    .B(_11392_),
    .Y(_11393_));
 a211o_1 _16400_ (.A1(net1153),
    .A2(_07073_),
    .B1(_07477_),
    .C1(_07550_),
    .X(_11394_));
 or2_1 _16401_ (.A(net715),
    .B(_10419_),
    .X(_11395_));
 and3b_1 _16402_ (.A_N(\digitop_pav2.sec_inst.ld_r.st[1] ),
    .B(\digitop_pav2.sec_inst.ld_r.st[0] ),
    .C(net716),
    .X(_11396_));
 nand3b_4 _16403_ (.A_N(\digitop_pav2.sec_inst.ld_r.st[1] ),
    .B(\digitop_pav2.sec_inst.ld_r.st[0] ),
    .C(net716),
    .Y(_11397_));
 nand2_1 _16404_ (.A(\digitop_pav2.sec_inst.shift_in.st[0] ),
    .B(\digitop_pav2.sec_inst.shift_in.st[1] ),
    .Y(_11398_));
 or2_1 _16405_ (.A(\digitop_pav2.sec_inst.shift_in.st[4] ),
    .B(_11398_),
    .X(_11399_));
 or2_2 _16406_ (.A(\digitop_pav2.sec_inst.shift_in.st[2] ),
    .B(\digitop_pav2.sec_inst.shift_in.st[3] ),
    .X(_11400_));
 or2_2 _16407_ (.A(_11399_),
    .B(_11400_),
    .X(_11401_));
 inv_2 _16408_ (.A(_11401_),
    .Y(_11402_));
 a21oi_1 _16409_ (.A1(\digitop_pav2.sec_inst.ld_r.st[0] ),
    .A2(\digitop_pav2.sec_inst.ld_r.st[1] ),
    .B1(net702),
    .Y(_11403_));
 a21o_1 _16410_ (.A1(\digitop_pav2.sec_inst.ld_r.st[0] ),
    .A2(\digitop_pav2.sec_inst.ld_r.st[1] ),
    .B1(net702),
    .X(_11404_));
 or2_1 _16411_ (.A(\digitop_pav2.sec_inst.ld_r.st[0] ),
    .B(\digitop_pav2.sec_inst.ld_r.st[1] ),
    .X(_11405_));
 a21bo_2 _16412_ (.A1(net702),
    .A2(_11405_),
    .B1_N(net717),
    .X(_11406_));
 nand2_2 _16413_ (.A(net716),
    .B(net682),
    .Y(_11407_));
 a31o_1 _16414_ (.A1(\digitop_pav2.sec_inst.shift_in.s4.q[0] ),
    .A2(net683),
    .A3(net577),
    .B1(_11407_),
    .X(_11408_));
 or3b_4 _16415_ (.A(\digitop_pav2.sec_inst.shift_in.st[4] ),
    .B(\digitop_pav2.sec_inst.shift_in.st[1] ),
    .C_N(\digitop_pav2.sec_inst.shift_in.st[0] ),
    .X(_11409_));
 nor2_1 _16416_ (.A(_11400_),
    .B(_11409_),
    .Y(_11410_));
 or2_1 _16417_ (.A(_11400_),
    .B(_11409_),
    .X(_11411_));
 and2_1 _16418_ (.A(net716),
    .B(_11405_),
    .X(_11412_));
 nand2_1 _16419_ (.A(net716),
    .B(\digitop_pav2.sec_inst.ld_r.st[1] ),
    .Y(_11413_));
 nor2_1 _16420_ (.A(\digitop_pav2.sec_inst.ld_r.st[0] ),
    .B(_11413_),
    .Y(_11414_));
 or2_1 _16421_ (.A(\digitop_pav2.sec_inst.ld_r.st[0] ),
    .B(_11413_),
    .X(_11415_));
 nand2_2 _16422_ (.A(_11397_),
    .B(net595),
    .Y(_11416_));
 nor2_2 _16423_ (.A(net683),
    .B(net598),
    .Y(_11417_));
 nand2b_2 _16424_ (.A_N(\digitop_pav2.sec_inst.shift_in.st[3] ),
    .B(\digitop_pav2.sec_inst.shift_in.st[2] ),
    .Y(_11418_));
 nor2_1 _16425_ (.A(_11409_),
    .B(_11418_),
    .Y(_11419_));
 or2_1 _16426_ (.A(_11409_),
    .B(_11418_),
    .X(_11420_));
 a31o_1 _16427_ (.A1(\digitop_pav2.sec_inst.shift_in.s6.q[0] ),
    .A2(net598),
    .A3(net594),
    .B1(_11408_),
    .X(_11421_));
 a31o_1 _16428_ (.A1(\digitop_pav2.sec_inst.shift_in.s2.q[0] ),
    .A2(_11411_),
    .A3(_11417_),
    .B1(_11421_),
    .X(_11422_));
 nand2b_2 _16429_ (.A_N(\digitop_pav2.sec_inst.shift_in.st[2] ),
    .B(\digitop_pav2.sec_inst.shift_in.st[3] ),
    .Y(_11423_));
 or2_4 _16430_ (.A(_11399_),
    .B(_11423_),
    .X(_11424_));
 inv_2 _16431_ (.A(_11424_),
    .Y(_11425_));
 nor2_2 _16432_ (.A(net596),
    .B(_11425_),
    .Y(_11426_));
 nor2_4 _16433_ (.A(_11409_),
    .B(_11423_),
    .Y(_11427_));
 nor2_2 _16434_ (.A(net598),
    .B(_11427_),
    .Y(_11428_));
 and3_1 _16435_ (.A(net702),
    .B(net716),
    .C(_11405_),
    .X(_11429_));
 nand2_1 _16436_ (.A(net702),
    .B(_11412_),
    .Y(_11430_));
 a221o_1 _16437_ (.A1(\digitop_pav2.sec_inst.shift_in.s12.q[0] ),
    .A2(_11426_),
    .B1(_11428_),
    .B2(\digitop_pav2.sec_inst.shift_in.s10.q[0] ),
    .C1(net575),
    .X(_11431_));
 nor2_1 _16438_ (.A(net682),
    .B(_11406_),
    .Y(_11432_));
 or2_2 _16439_ (.A(net682),
    .B(_11406_),
    .X(_11433_));
 or2_2 _16440_ (.A(_11399_),
    .B(_11418_),
    .X(_11434_));
 inv_2 _16441_ (.A(net574),
    .Y(_11435_));
 a21o_1 _16442_ (.A1(\digitop_pav2.sec_inst.shift_in.s8.q[0] ),
    .A2(net574),
    .B1(_11433_),
    .X(_11436_));
 o211a_1 _16443_ (.A1(net1135),
    .A2(net717),
    .B1(net601),
    .C1(_11436_),
    .X(_11437_));
 a32o_1 _16444_ (.A1(_11422_),
    .A2(_11431_),
    .A3(_11437_),
    .B1(net602),
    .B2(_08877_),
    .X(_11438_));
 nand2_1 _16445_ (.A(net535),
    .B(_11438_),
    .Y(_11439_));
 a21oi_2 _16446_ (.A1(_11394_),
    .A2(_11439_),
    .B1(_07520_),
    .Y(_11440_));
 nor2_8 _16447_ (.A(net471),
    .B(_11223_),
    .Y(_11441_));
 or2_1 _16448_ (.A(net471),
    .B(_11223_),
    .X(_11442_));
 nor2_1 _16449_ (.A(net187),
    .B(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_9.Y ),
    .Y(_11443_));
 nand2_2 _16450_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_9.Y ),
    .B(net183),
    .Y(_11444_));
 nor2_4 _16451_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_9.Y ),
    .B(net183),
    .Y(_11445_));
 nand2_2 _16452_ (.A(net187),
    .B(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_9.Y ),
    .Y(_11446_));
 nor2_1 _16453_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_9.Y ),
    .B(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_9.Y ),
    .Y(_11447_));
 or2_1 _16454_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_9.Y ),
    .B(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_9.Y ),
    .X(_11448_));
 a221o_1 _16455_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[8] ),
    .A2(net184),
    .B1(net165),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[8] ),
    .C1(net178),
    .X(_11449_));
 a21o_1 _16456_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[8] ),
    .A2(net169),
    .B1(_11449_),
    .X(_11450_));
 o21ai_2 _16457_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[8] ),
    .A2(net172),
    .B1(_11450_),
    .Y(_11451_));
 nor2_1 _16458_ (.A(net347),
    .B(_11451_),
    .Y(_11452_));
 a221o_1 _16459_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[15] ),
    .A2(net184),
    .B1(net166),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[15] ),
    .C1(net176),
    .X(_11453_));
 a21o_1 _16460_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[15] ),
    .A2(net162),
    .B1(_11453_),
    .X(_11454_));
 o21ai_1 _16461_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[15] ),
    .A2(net172),
    .B1(_11454_),
    .Y(_11455_));
 or2_4 _16462_ (.A(net347),
    .B(_11455_),
    .X(_11456_));
 inv_2 _16463_ (.A(_11456_),
    .Y(_11457_));
 a22o_1 _16464_ (.A1(_11452_),
    .A2(_11455_),
    .B1(_11457_),
    .B2(_11451_),
    .X(_11458_));
 a221o_1 _16465_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[7] ),
    .A2(net184),
    .B1(net162),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ),
    .C1(net176),
    .X(_11459_));
 a21o_1 _16466_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[7] ),
    .A2(net166),
    .B1(_11459_),
    .X(_11460_));
 o21ai_4 _16467_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ),
    .A2(net172),
    .B1(_11460_),
    .Y(_11461_));
 nor2_2 _16468_ (.A(net348),
    .B(_11461_),
    .Y(_11462_));
 or2_2 _16469_ (.A(net348),
    .B(_11461_),
    .X(_11463_));
 a221o_1 _16470_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[0] ),
    .A2(net185),
    .B1(net167),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[0] ),
    .C1(net177),
    .X(_11464_));
 a21o_1 _16471_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[0] ),
    .A2(net163),
    .B1(_11464_),
    .X(_11465_));
 o21ai_2 _16472_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[0] ),
    .A2(net174),
    .B1(_11465_),
    .Y(_11466_));
 nor2_2 _16473_ (.A(net347),
    .B(_11466_),
    .Y(_11467_));
 a221o_1 _16474_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[8] ),
    .A2(net184),
    .B1(net162),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[8] ),
    .C1(net176),
    .X(_11468_));
 a21o_1 _16475_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[8] ),
    .A2(net169),
    .B1(_11468_),
    .X(_11469_));
 o21ai_2 _16476_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[8] ),
    .A2(net173),
    .B1(_11469_),
    .Y(_11470_));
 nor2_1 _16477_ (.A(net347),
    .B(_11470_),
    .Y(_11471_));
 a22o_1 _16478_ (.A1(_11467_),
    .A2(_11470_),
    .B1(_11471_),
    .B2(_11466_),
    .X(_11472_));
 xnor2_1 _16479_ (.A(_11463_),
    .B(_11472_),
    .Y(_11473_));
 nand2_1 _16480_ (.A(_11458_),
    .B(_11473_),
    .Y(_11474_));
 or2_1 _16481_ (.A(_11458_),
    .B(_11473_),
    .X(_11475_));
 a31o_1 _16482_ (.A1(net467),
    .A2(_11474_),
    .A3(_11475_),
    .B1(_11440_),
    .X(_11476_));
 or2_1 _16483_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[0] ),
    .X(_11477_));
 nand2_1 _16484_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[0] ),
    .Y(_11478_));
 o21ai_1 _16485_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[0] ),
    .B1(net434),
    .Y(_11479_));
 a21oi_1 _16486_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[0] ),
    .B1(_11479_),
    .Y(_11480_));
 a31o_1 _16487_ (.A1(net420),
    .A2(_11477_),
    .A3(_11478_),
    .B1(_11480_),
    .X(_11481_));
 or4b_1 _16488_ (.A(_11393_),
    .B(_11476_),
    .C(_11481_),
    .D_N(net161),
    .X(_11482_));
 xnor2_1 _16489_ (.A(_11452_),
    .B(_11456_),
    .Y(_11483_));
 o21a_1 _16490_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[0] ),
    .A2(net161),
    .B1(_11482_),
    .X(_00357_));
 nand2_1 _16491_ (.A(net237),
    .B(_11281_),
    .Y(_11484_));
 o31a_1 _16492_ (.A1(net237),
    .A2(_11261_),
    .A3(_11348_),
    .B1(_11484_),
    .X(_11485_));
 nand2_1 _16493_ (.A(_11288_),
    .B(_11295_),
    .Y(_11486_));
 and3_1 _16494_ (.A(net237),
    .B(_11292_),
    .C(_11486_),
    .X(_11487_));
 or3_1 _16495_ (.A(net223),
    .B(_11307_),
    .C(_11373_),
    .X(_11488_));
 a21oi_1 _16496_ (.A1(_11315_),
    .A2(_11329_),
    .B1(_11317_),
    .Y(_11489_));
 nor2_1 _16497_ (.A(_11275_),
    .B(_11368_),
    .Y(_11490_));
 o221a_1 _16498_ (.A1(_11261_),
    .A2(_11312_),
    .B1(_11368_),
    .B2(_11275_),
    .C1(net229),
    .X(_11491_));
 nand2_1 _16499_ (.A(_11264_),
    .B(_11294_),
    .Y(_11492_));
 a221o_1 _16500_ (.A1(_11290_),
    .A2(_11372_),
    .B1(_11492_),
    .B2(_11342_),
    .C1(net229),
    .X(_11493_));
 nand2_1 _16501_ (.A(net240),
    .B(_11339_),
    .Y(_11494_));
 nor2_2 _16502_ (.A(net288),
    .B(net200),
    .Y(_11495_));
 or2_1 _16503_ (.A(net237),
    .B(_11495_),
    .X(_11496_));
 o32a_1 _16504_ (.A1(_11276_),
    .A2(_11338_),
    .A3(_11496_),
    .B1(_11494_),
    .B2(_11287_),
    .X(_11497_));
 o21ai_1 _16505_ (.A1(net222),
    .A2(_11497_),
    .B1(_11493_),
    .Y(_11498_));
 nor2_1 _16506_ (.A(_11320_),
    .B(_11372_),
    .Y(_02152_));
 o211a_1 _16507_ (.A1(net238),
    .A2(_11340_),
    .B1(_02152_),
    .C1(net222),
    .X(_02153_));
 o221a_1 _16508_ (.A1(net227),
    .A2(_11485_),
    .B1(_11487_),
    .B2(_11488_),
    .C1(net284),
    .X(_02154_));
 a211oi_1 _16509_ (.A1(net282),
    .A2(_11498_),
    .B1(_02154_),
    .C1(net248),
    .Y(_02155_));
 a41o_1 _16510_ (.A1(_11264_),
    .A2(net227),
    .A3(_11316_),
    .A4(_11380_),
    .B1(net284),
    .X(_02156_));
 o32a_1 _16511_ (.A1(net282),
    .A2(_11489_),
    .A3(_11491_),
    .B1(_02153_),
    .B2(_02156_),
    .X(_02157_));
 a211o_1 _16512_ (.A1(net248),
    .A2(_02157_),
    .B1(_02155_),
    .C1(_11357_),
    .X(_02158_));
 and2_1 _16513_ (.A(net245),
    .B(net236),
    .X(_02159_));
 nand2_2 _16514_ (.A(net242),
    .B(net235),
    .Y(_02160_));
 o221a_1 _16515_ (.A1(net243),
    .A2(_11486_),
    .B1(_02160_),
    .B2(_11280_),
    .C1(net248),
    .X(_02161_));
 o221a_1 _16516_ (.A1(_11289_),
    .A2(_11329_),
    .B1(_11484_),
    .B2(_11251_),
    .C1(net251),
    .X(_02162_));
 nor2_1 _16517_ (.A(_11282_),
    .B(_11340_),
    .Y(_02163_));
 or2_1 _16518_ (.A(_11338_),
    .B(_11367_),
    .X(_02164_));
 nor2_1 _16519_ (.A(net237),
    .B(_02163_),
    .Y(_02165_));
 a211o_1 _16520_ (.A1(net251),
    .A2(_11311_),
    .B1(_02165_),
    .C1(net224),
    .X(_02166_));
 o311a_1 _16521_ (.A1(net228),
    .A2(_02161_),
    .A3(_02162_),
    .B1(_02166_),
    .C1(net284),
    .X(_02167_));
 a21o_1 _16522_ (.A1(_11380_),
    .A2(_02160_),
    .B1(_11495_),
    .X(_02168_));
 nor2_1 _16523_ (.A(_11276_),
    .B(_11312_),
    .Y(_02169_));
 nor2_1 _16524_ (.A(net289),
    .B(_11262_),
    .Y(_02170_));
 nor2_1 _16525_ (.A(_11289_),
    .B(_11363_),
    .Y(_02171_));
 nand2_1 _16526_ (.A(_11252_),
    .B(_02169_),
    .Y(_02172_));
 nand2_1 _16527_ (.A(net242),
    .B(_11363_),
    .Y(_02173_));
 and4bb_1 _16528_ (.A_N(net251),
    .B_N(_11495_),
    .C(_02172_),
    .D(_02173_),
    .X(_02174_));
 a311o_1 _16529_ (.A1(net251),
    .A2(_11316_),
    .A3(_02168_),
    .B1(_02174_),
    .C1(net227),
    .X(_02175_));
 or3_1 _16530_ (.A(net237),
    .B(_11261_),
    .C(_11340_),
    .X(_02176_));
 o211a_1 _16531_ (.A1(net243),
    .A2(_11310_),
    .B1(_02176_),
    .C1(net251),
    .X(_02177_));
 nor2_1 _16532_ (.A(_11276_),
    .B(_11495_),
    .Y(_02178_));
 a311o_1 _16533_ (.A1(net248),
    .A2(_11321_),
    .A3(_02178_),
    .B1(_02177_),
    .C1(net224),
    .X(_02179_));
 a31o_1 _16534_ (.A1(net282),
    .A2(_02175_),
    .A3(_02179_),
    .B1(_02167_),
    .X(_02180_));
 o211a_2 _16535_ (.A1(net280),
    .A2(_02180_),
    .B1(_02158_),
    .C1(_11361_),
    .X(_02181_));
 and2_2 _16536_ (.A(net472),
    .B(_02181_),
    .X(_02182_));
 a211o_1 _16537_ (.A1(net1153),
    .A2(net1132),
    .B1(_07477_),
    .C1(net1017),
    .X(_02183_));
 a31o_1 _16538_ (.A1(\digitop_pav2.sec_inst.shift_in.s2.q[1] ),
    .A2(net599),
    .A3(_11417_),
    .B1(_11407_),
    .X(_02184_));
 a31o_1 _16539_ (.A1(\digitop_pav2.sec_inst.shift_in.s6.q[1] ),
    .A2(net598),
    .A3(net594),
    .B1(_02184_),
    .X(_02185_));
 a31o_1 _16540_ (.A1(\digitop_pav2.sec_inst.shift_in.s4.q[1] ),
    .A2(net683),
    .A3(_11401_),
    .B1(_02185_),
    .X(_02186_));
 a221o_1 _16541_ (.A1(\digitop_pav2.sec_inst.shift_in.s12.q[1] ),
    .A2(_11426_),
    .B1(_11428_),
    .B2(\digitop_pav2.sec_inst.shift_in.s10.q[1] ),
    .C1(net575),
    .X(_02187_));
 a21o_1 _16542_ (.A1(\digitop_pav2.sec_inst.shift_in.s8.q[1] ),
    .A2(net574),
    .B1(_11433_),
    .X(_02188_));
 o211a_1 _16543_ (.A1(net1132),
    .A2(net717),
    .B1(net601),
    .C1(_02188_),
    .X(_02189_));
 a32o_1 _16544_ (.A1(_02186_),
    .A2(_02187_),
    .A3(_02189_),
    .B1(net602),
    .B2(_08889_),
    .X(_02190_));
 a22o_1 _16545_ (.A1(net1255),
    .A2(_02183_),
    .B1(_02190_),
    .B2(net534),
    .X(_02191_));
 and2_2 _16546_ (.A(net398),
    .B(_02191_),
    .X(_02192_));
 a22o_1 _16547_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[9] ),
    .A2(net162),
    .B1(_11445_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[9] ),
    .X(_02193_));
 a211o_1 _16548_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[9] ),
    .A2(net166),
    .B1(net176),
    .C1(_02193_),
    .X(_02194_));
 o21ai_1 _16549_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[9] ),
    .A2(net172),
    .B1(_02194_),
    .Y(_02195_));
 or2_2 _16550_ (.A(net347),
    .B(_02195_),
    .X(_02196_));
 inv_2 _16551_ (.A(_02196_),
    .Y(_02197_));
 a221o_1 _16552_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[1] ),
    .A2(net185),
    .B1(net163),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[1] ),
    .C1(net177),
    .X(_02198_));
 a21o_1 _16553_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[1] ),
    .A2(net167),
    .B1(_02198_),
    .X(_02199_));
 o21ai_2 _16554_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[1] ),
    .A2(net174),
    .B1(_02199_),
    .Y(_02200_));
 or2_2 _16555_ (.A(net347),
    .B(_02200_),
    .X(_02201_));
 inv_2 _16556_ (.A(_02201_),
    .Y(_02202_));
 mux2_1 _16557_ (.A0(_02200_),
    .A1(_02202_),
    .S(_02196_),
    .X(_02203_));
 a221o_1 _16558_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[0] ),
    .A2(net185),
    .B1(net163),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ),
    .C1(net177),
    .X(_02204_));
 a21o_1 _16559_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[0] ),
    .A2(net167),
    .B1(_02204_),
    .X(_02205_));
 o21ai_2 _16560_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[0] ),
    .A2(net174),
    .B1(_02205_),
    .Y(_02206_));
 nor2_2 _16561_ (.A(net347),
    .B(_02206_),
    .Y(_02207_));
 a22o_1 _16562_ (.A1(_11462_),
    .A2(_02206_),
    .B1(_02207_),
    .B2(_11461_),
    .X(_02208_));
 a22o_1 _16563_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[9] ),
    .A2(net162),
    .B1(_11445_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[9] ),
    .X(_02209_));
 a211o_1 _16564_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[9] ),
    .A2(net166),
    .B1(net176),
    .C1(_02209_),
    .X(_02210_));
 o21ai_1 _16565_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[9] ),
    .A2(net172),
    .B1(_02210_),
    .Y(_02211_));
 or2_2 _16566_ (.A(net347),
    .B(_02211_),
    .X(_02212_));
 inv_2 _16567_ (.A(_02212_),
    .Y(_02213_));
 o21ai_1 _16568_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[1] ),
    .B1(net432),
    .Y(_02214_));
 a21oi_1 _16569_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[1] ),
    .B1(_02214_),
    .Y(_02215_));
 or2_1 _16570_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[1] ),
    .X(_02216_));
 nand2_1 _16571_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[1] ),
    .Y(_02217_));
 a31o_1 _16572_ (.A1(net418),
    .A2(_02216_),
    .A3(_02217_),
    .B1(_02215_),
    .X(_02218_));
 xnor2_2 _16573_ (.A(_11463_),
    .B(_02207_),
    .Y(_02219_));
 xnor2_1 _16574_ (.A(_02203_),
    .B(_02219_),
    .Y(_02220_));
 xnor2_1 _16575_ (.A(_11483_),
    .B(_02213_),
    .Y(_02221_));
 nor2_1 _16576_ (.A(_02220_),
    .B(_02221_),
    .Y(_02222_));
 nand2_1 _16577_ (.A(_02220_),
    .B(_02221_),
    .Y(_02223_));
 and3b_1 _16578_ (.A_N(_02222_),
    .B(_02223_),
    .C(net466),
    .X(_02224_));
 or4_1 _16579_ (.A(_02182_),
    .B(_02192_),
    .C(_02218_),
    .D(_02224_),
    .X(_02225_));
 mux2_1 _16580_ (.A0(\digitop_pav2.aes128_inst.aes128_regs.state2_r[1] ),
    .A1(_02225_),
    .S(net161),
    .X(_00358_));
 o21ba_1 _16581_ (.A1(_11341_),
    .A2(_02170_),
    .B1_N(_11370_),
    .X(_02226_));
 or3b_1 _16582_ (.A(_11347_),
    .B(net241),
    .C_N(net200),
    .X(_02227_));
 nor2_1 _16583_ (.A(_11264_),
    .B(_11294_),
    .Y(_02228_));
 a211o_1 _16584_ (.A1(_02178_),
    .A2(_02227_),
    .B1(_02228_),
    .C1(net229),
    .X(_02229_));
 o211a_1 _16585_ (.A1(net223),
    .A2(_02226_),
    .B1(_02229_),
    .C1(net286),
    .X(_02230_));
 nand2_1 _16586_ (.A(_11296_),
    .B(_11310_),
    .Y(_02231_));
 nor2_1 _16587_ (.A(net239),
    .B(_11281_),
    .Y(_02232_));
 nand2_1 _16588_ (.A(net230),
    .B(_02160_),
    .Y(_02233_));
 a211o_1 _16589_ (.A1(net239),
    .A2(_02231_),
    .B1(_02232_),
    .C1(_02233_),
    .X(_02234_));
 o211a_1 _16590_ (.A1(net238),
    .A2(_11290_),
    .B1(_02160_),
    .C1(net223),
    .X(_02235_));
 nand2_1 _16591_ (.A(net240),
    .B(_11278_),
    .Y(_02236_));
 o21ai_1 _16592_ (.A1(_11289_),
    .A2(_02236_),
    .B1(_02235_),
    .Y(_02237_));
 a31o_1 _16593_ (.A1(net241),
    .A2(_11308_),
    .A3(_11364_),
    .B1(net226),
    .X(_02238_));
 o21ai_2 _16594_ (.A1(_11338_),
    .A2(_11380_),
    .B1(_11346_),
    .Y(_02239_));
 a31o_1 _16595_ (.A1(net241),
    .A2(net288),
    .A3(_11262_),
    .B1(net232),
    .X(_02240_));
 o221a_1 _16596_ (.A1(_11381_),
    .A2(_02238_),
    .B1(_02239_),
    .B2(_02240_),
    .C1(net285),
    .X(_02241_));
 o32a_1 _16597_ (.A1(_11261_),
    .A2(_11287_),
    .A3(_11312_),
    .B1(_11348_),
    .B2(_11264_),
    .X(_02242_));
 nand2_1 _16598_ (.A(net225),
    .B(_02242_),
    .Y(_02243_));
 a221o_1 _16599_ (.A1(net237),
    .A2(_11295_),
    .B1(_11363_),
    .B2(_11379_),
    .C1(net225),
    .X(_02244_));
 a21oi_1 _16600_ (.A1(_02243_),
    .A2(_02244_),
    .B1(net285),
    .Y(_02245_));
 a31o_1 _16601_ (.A1(net246),
    .A2(_11242_),
    .A3(_11262_),
    .B1(net232),
    .X(_02246_));
 a21o_1 _16602_ (.A1(net241),
    .A2(_11297_),
    .B1(_02246_),
    .X(_02247_));
 or2_1 _16603_ (.A(_11275_),
    .B(_11484_),
    .X(_02248_));
 or3b_1 _16604_ (.A(net223),
    .B(_11307_),
    .C_N(_02248_),
    .X(_02249_));
 a221o_1 _16605_ (.A1(net240),
    .A2(_11293_),
    .B1(_02159_),
    .B2(_11280_),
    .C1(net225),
    .X(_02250_));
 o211a_1 _16606_ (.A1(_11369_),
    .A2(_02240_),
    .B1(_02250_),
    .C1(net285),
    .X(_02251_));
 a31o_1 _16607_ (.A1(net240),
    .A2(_11364_),
    .A3(_11386_),
    .B1(_11379_),
    .X(_02252_));
 nand2_1 _16608_ (.A(net233),
    .B(_02252_),
    .Y(_02253_));
 a211o_1 _16609_ (.A1(_11288_),
    .A2(_11311_),
    .B1(_11381_),
    .C1(net233),
    .X(_02254_));
 nand2_1 _16610_ (.A(_11277_),
    .B(_11379_),
    .Y(_02255_));
 o21a_1 _16611_ (.A1(_11251_),
    .A2(_02236_),
    .B1(_02255_),
    .X(_02256_));
 a31o_1 _16612_ (.A1(net240),
    .A2(_11277_),
    .A3(_11339_),
    .B1(net233),
    .X(_02257_));
 o221a_1 _16613_ (.A1(net225),
    .A2(_02256_),
    .B1(_02257_),
    .B2(_02165_),
    .C1(net285),
    .X(_02258_));
 a311o_1 _16614_ (.A1(net283),
    .A2(_02247_),
    .A3(_02249_),
    .B1(_02251_),
    .C1(_11357_),
    .X(_02259_));
 o311a_1 _16615_ (.A1(net280),
    .A2(_02241_),
    .A3(_02245_),
    .B1(_02259_),
    .C1(net252),
    .X(_02260_));
 a31o_1 _16616_ (.A1(net283),
    .A2(_02253_),
    .A3(_02254_),
    .B1(_02258_),
    .X(_02261_));
 nand2_1 _16617_ (.A(net280),
    .B(_02261_),
    .Y(_02262_));
 a311o_1 _16618_ (.A1(net282),
    .A2(_02234_),
    .A3(_02237_),
    .B1(net280),
    .C1(_02230_),
    .X(_02263_));
 a31o_2 _16619_ (.A1(net249),
    .A2(_02262_),
    .A3(_02263_),
    .B1(_02260_),
    .X(_02264_));
 nor2_2 _16620_ (.A(_07092_),
    .B(_02264_),
    .Y(_02265_));
 o21ai_1 _16621_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[2] ),
    .B1(net435),
    .Y(_02266_));
 a21oi_1 _16622_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[2] ),
    .B1(_02266_),
    .Y(_02267_));
 a21boi_1 _16623_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[2] ),
    .B1_N(net421),
    .Y(_02268_));
 o21a_1 _16624_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[2] ),
    .B1(_02268_),
    .X(_02269_));
 a21oi_2 _16625_ (.A1(_07025_),
    .A2(net1049),
    .B1(net1155),
    .Y(_02270_));
 a211o_1 _16626_ (.A1(net1153),
    .A2(net1130),
    .B1(net1017),
    .C1(_02270_),
    .X(_02271_));
 a31o_1 _16627_ (.A1(\digitop_pav2.sec_inst.shift_in.s2.q[2] ),
    .A2(net599),
    .A3(_11417_),
    .B1(_11407_),
    .X(_02272_));
 a31o_1 _16628_ (.A1(\digitop_pav2.sec_inst.shift_in.s6.q[2] ),
    .A2(net598),
    .A3(net594),
    .B1(_02272_),
    .X(_02273_));
 a31o_1 _16629_ (.A1(\digitop_pav2.sec_inst.shift_in.s4.q[2] ),
    .A2(net683),
    .A3(_11401_),
    .B1(_02273_),
    .X(_02274_));
 a221o_1 _16630_ (.A1(\digitop_pav2.sec_inst.shift_in.s12.q[2] ),
    .A2(_11426_),
    .B1(_11428_),
    .B2(\digitop_pav2.sec_inst.shift_in.s10.q[2] ),
    .C1(net576),
    .X(_02275_));
 a21o_1 _16631_ (.A1(\digitop_pav2.sec_inst.shift_in.s8.q[2] ),
    .A2(net574),
    .B1(_11433_),
    .X(_02276_));
 o211a_1 _16632_ (.A1(net1130),
    .A2(net717),
    .B1(net601),
    .C1(_02276_),
    .X(_02277_));
 a32o_1 _16633_ (.A1(_02274_),
    .A2(_02275_),
    .A3(_02277_),
    .B1(net603),
    .B2(_08891_),
    .X(_02278_));
 a22o_1 _16634_ (.A1(net1255),
    .A2(_02271_),
    .B1(_02278_),
    .B2(net534),
    .X(_02279_));
 and2_2 _16635_ (.A(_07519_),
    .B(_02279_),
    .X(_02280_));
 a221o_1 _16636_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[10] ),
    .A2(net184),
    .B1(net166),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[10] ),
    .C1(net176),
    .X(_02281_));
 a21o_1 _16637_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[10] ),
    .A2(net162),
    .B1(_02281_),
    .X(_02282_));
 o21ai_1 _16638_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[10] ),
    .A2(net172),
    .B1(_02282_),
    .Y(_02283_));
 or2_2 _16639_ (.A(net348),
    .B(_02283_),
    .X(_02284_));
 inv_2 _16640_ (.A(_02284_),
    .Y(_02285_));
 a22o_1 _16641_ (.A1(_02213_),
    .A2(_02283_),
    .B1(_02285_),
    .B2(_02211_),
    .X(_02286_));
 a221o_1 _16642_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[1] ),
    .A2(net185),
    .B1(net167),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[1] ),
    .C1(net177),
    .X(_02287_));
 a21o_1 _16643_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[1] ),
    .A2(net163),
    .B1(_02287_),
    .X(_02288_));
 o21ai_1 _16644_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[1] ),
    .A2(net174),
    .B1(_02288_),
    .Y(_02289_));
 or2_1 _16645_ (.A(net347),
    .B(_02289_),
    .X(_02290_));
 inv_2 _16646_ (.A(_02290_),
    .Y(_02291_));
 a22o_1 _16647_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[2] ),
    .A2(net185),
    .B1(net183),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[2] ),
    .X(_02292_));
 a211o_1 _16648_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[2] ),
    .A2(net167),
    .B1(net177),
    .C1(_02292_),
    .X(_02293_));
 o21ai_2 _16649_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[2] ),
    .A2(net174),
    .B1(_02293_),
    .Y(_02294_));
 nor2_2 _16650_ (.A(net347),
    .B(_02294_),
    .Y(_02295_));
 a221o_1 _16651_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[10] ),
    .A2(net184),
    .B1(net162),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ),
    .C1(net176),
    .X(_02296_));
 a21o_1 _16652_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ),
    .A2(net166),
    .B1(_02296_),
    .X(_02297_));
 o21ai_1 _16653_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[10] ),
    .A2(net172),
    .B1(_02297_),
    .Y(_02298_));
 or2_2 _16654_ (.A(net348),
    .B(_02298_),
    .X(_02299_));
 xor2_1 _16655_ (.A(_02295_),
    .B(_02299_),
    .X(_02300_));
 xnor2_1 _16656_ (.A(_02291_),
    .B(_02300_),
    .Y(_02301_));
 nor2_1 _16657_ (.A(_02286_),
    .B(_02301_),
    .Y(_02302_));
 nand2_1 _16658_ (.A(_02286_),
    .B(_02301_),
    .Y(_02303_));
 and3b_1 _16659_ (.A_N(_02302_),
    .B(_02303_),
    .C(net466),
    .X(_02304_));
 or2_1 _16660_ (.A(_02280_),
    .B(_02304_),
    .X(_02305_));
 or4b_1 _16661_ (.A(_02267_),
    .B(_02269_),
    .C(_02305_),
    .D_N(net161),
    .X(_02306_));
 o22a_1 _16662_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[2] ),
    .A2(net161),
    .B1(_02265_),
    .B2(_02306_),
    .X(_00359_));
 o22a_1 _16663_ (.A1(net245),
    .A2(_11285_),
    .B1(_11289_),
    .B2(_11329_),
    .X(_02307_));
 nor2_1 _16664_ (.A(net233),
    .B(_02307_),
    .Y(_02308_));
 o211a_1 _16665_ (.A1(_11334_),
    .A2(_02236_),
    .B1(_02173_),
    .C1(net233),
    .X(_02309_));
 nand2_1 _16666_ (.A(net244),
    .B(_11310_),
    .Y(_02310_));
 inv_2 _16667_ (.A(_02310_),
    .Y(_02311_));
 o211a_1 _16668_ (.A1(_11291_),
    .A2(_02310_),
    .B1(_02152_),
    .C1(net223),
    .X(_02312_));
 a311o_1 _16669_ (.A1(net228),
    .A2(_11364_),
    .A3(_02173_),
    .B1(_02312_),
    .C1(net284),
    .X(_02313_));
 o311a_1 _16670_ (.A1(net282),
    .A2(_02308_),
    .A3(_02309_),
    .B1(_02313_),
    .C1(net280),
    .X(_02314_));
 nand2_1 _16671_ (.A(net242),
    .B(_11315_),
    .Y(_02315_));
 o311a_1 _16672_ (.A1(net242),
    .A2(_11287_),
    .A3(_02170_),
    .B1(_02315_),
    .C1(net228),
    .X(_02316_));
 a21oi_1 _16673_ (.A1(net237),
    .A2(_11363_),
    .B1(net227),
    .Y(_02317_));
 a311o_1 _16674_ (.A1(_11292_),
    .A2(_11294_),
    .A3(_02317_),
    .B1(_02316_),
    .C1(net282),
    .X(_02318_));
 a21oi_2 _16675_ (.A1(_11288_),
    .A2(_11292_),
    .B1(net245),
    .Y(_02319_));
 o21a_1 _16676_ (.A1(_02165_),
    .A2(_02319_),
    .B1(net233),
    .X(_02320_));
 o311a_1 _16677_ (.A1(net284),
    .A2(_02235_),
    .A3(_02320_),
    .B1(_02318_),
    .C1(_11357_),
    .X(_02321_));
 a21oi_1 _16678_ (.A1(net200),
    .A2(_11284_),
    .B1(net240),
    .Y(_02322_));
 o21ai_1 _16679_ (.A1(_11263_),
    .A2(_02322_),
    .B1(net226),
    .Y(_02323_));
 a32o_1 _16680_ (.A1(net239),
    .A2(_11294_),
    .A3(_11363_),
    .B1(_11330_),
    .B2(_11283_),
    .X(_02324_));
 and3_1 _16681_ (.A(net237),
    .B(_11278_),
    .C(net200),
    .X(_02325_));
 a2111o_1 _16682_ (.A1(net244),
    .A2(_11315_),
    .B1(_02325_),
    .C1(net229),
    .D1(_11307_),
    .X(_02326_));
 a21oi_1 _16683_ (.A1(net243),
    .A2(_02171_),
    .B1(net224),
    .Y(_02327_));
 a31o_1 _16684_ (.A1(_11262_),
    .A2(_11288_),
    .A3(_11320_),
    .B1(net229),
    .X(_02328_));
 a31o_1 _16685_ (.A1(_11278_),
    .A2(net200),
    .A3(_11321_),
    .B1(_02328_),
    .X(_02329_));
 a21bo_1 _16686_ (.A1(_11486_),
    .A2(_02327_),
    .B1_N(_02329_),
    .X(_02330_));
 a211o_1 _16687_ (.A1(net238),
    .A2(_11331_),
    .B1(_02311_),
    .C1(net230),
    .X(_02331_));
 or3b_1 _16688_ (.A(_02232_),
    .B(_02233_),
    .C_N(_02236_),
    .X(_02332_));
 o211a_1 _16689_ (.A1(net224),
    .A2(_02324_),
    .B1(_02323_),
    .C1(net282),
    .X(_02333_));
 a211oi_1 _16690_ (.A1(net284),
    .A2(_02330_),
    .B1(_02333_),
    .C1(_11357_),
    .Y(_02334_));
 o311a_1 _16691_ (.A1(net222),
    .A2(_11372_),
    .A3(_11490_),
    .B1(_02326_),
    .C1(net282),
    .X(_02335_));
 a311o_1 _16692_ (.A1(net286),
    .A2(_02331_),
    .A3(_02332_),
    .B1(_02335_),
    .C1(net280),
    .X(_02336_));
 nand2_1 _16693_ (.A(net250),
    .B(_02336_),
    .Y(_02337_));
 o32a_4 _16694_ (.A1(net248),
    .A2(_02314_),
    .A3(_02321_),
    .B1(_02334_),
    .B2(_02337_),
    .X(_02338_));
 and2_2 _16695_ (.A(net472),
    .B(_02338_),
    .X(_02339_));
 o21ai_1 _16696_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[3] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[3] ),
    .B1(net436),
    .Y(_02340_));
 a21oi_1 _16697_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[3] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[3] ),
    .B1(_02340_),
    .Y(_02341_));
 or2_1 _16698_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[3] ),
    .X(_02342_));
 nand2_1 _16699_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[3] ),
    .Y(_02343_));
 a31o_1 _16700_ (.A1(net422),
    .A2(_02342_),
    .A3(_02343_),
    .B1(_02341_),
    .X(_02344_));
 a211o_1 _16701_ (.A1(net1153),
    .A2(net1126),
    .B1(_07477_),
    .C1(net1017),
    .X(_02345_));
 a31o_1 _16702_ (.A1(\digitop_pav2.sec_inst.shift_in.s4.q[3] ),
    .A2(net683),
    .A3(net577),
    .B1(_11407_),
    .X(_02346_));
 a31o_1 _16703_ (.A1(\digitop_pav2.sec_inst.shift_in.s6.q[3] ),
    .A2(net598),
    .A3(net594),
    .B1(_02346_),
    .X(_02347_));
 a31o_1 _16704_ (.A1(\digitop_pav2.sec_inst.shift_in.s2.q[3] ),
    .A2(net599),
    .A3(_11417_),
    .B1(_02347_),
    .X(_02348_));
 a221o_1 _16705_ (.A1(\digitop_pav2.sec_inst.shift_in.s12.q[3] ),
    .A2(_11426_),
    .B1(_11428_),
    .B2(\digitop_pav2.sec_inst.shift_in.s10.q[3] ),
    .C1(net576),
    .X(_02349_));
 a21o_1 _16706_ (.A1(\digitop_pav2.sec_inst.shift_in.s8.q[3] ),
    .A2(net574),
    .B1(_11433_),
    .X(_02350_));
 o211a_1 _16707_ (.A1(net1126),
    .A2(net717),
    .B1(net601),
    .C1(_02350_),
    .X(_02351_));
 a32o_1 _16708_ (.A1(_02348_),
    .A2(_02349_),
    .A3(_02351_),
    .B1(net602),
    .B2(_08886_),
    .X(_02352_));
 a22o_1 _16709_ (.A1(net1255),
    .A2(_02345_),
    .B1(_02352_),
    .B2(net534),
    .X(_02353_));
 and2_2 _16710_ (.A(net398),
    .B(_02353_),
    .X(_02354_));
 a22o_1 _16711_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[2] ),
    .A2(net163),
    .B1(_11445_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[2] ),
    .X(_02355_));
 a211o_1 _16712_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[2] ),
    .A2(net167),
    .B1(net177),
    .C1(_02355_),
    .X(_02356_));
 o211ai_4 _16713_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ),
    .A2(net174),
    .B1(_02356_),
    .C1(_11441_),
    .Y(_02357_));
 mux2_1 _16714_ (.A0(_11461_),
    .A1(_11462_),
    .S(_02357_),
    .X(_02358_));
 a221o_1 _16715_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[3] ),
    .A2(net185),
    .B1(net167),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[3] ),
    .C1(net177),
    .X(_02359_));
 a21o_1 _16716_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[3] ),
    .A2(net163),
    .B1(_02359_),
    .X(_02360_));
 o21ai_1 _16717_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[3] ),
    .A2(net174),
    .B1(_02360_),
    .Y(_02361_));
 or2_2 _16718_ (.A(net348),
    .B(_02361_),
    .X(_02362_));
 inv_2 _16719_ (.A(_02362_),
    .Y(_02363_));
 a221o_1 _16720_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[11] ),
    .A2(net184),
    .B1(net169),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[11] ),
    .C1(net176),
    .X(_02364_));
 a21o_1 _16721_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[11] ),
    .A2(net165),
    .B1(_02364_),
    .X(_02365_));
 o21ai_1 _16722_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[11] ),
    .A2(net173),
    .B1(_02365_),
    .Y(_02366_));
 inv_2 _16723_ (.A(_02366_),
    .Y(_02367_));
 or2_1 _16724_ (.A(net349),
    .B(_02366_),
    .X(_02368_));
 a22o_1 _16725_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[11] ),
    .A2(net165),
    .B1(_11445_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[11] ),
    .X(_02369_));
 a211o_1 _16726_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[11] ),
    .A2(net166),
    .B1(net178),
    .C1(_02369_),
    .X(_02370_));
 o21ai_1 _16727_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[11] ),
    .A2(net173),
    .B1(_02370_),
    .Y(_02371_));
 or2_2 _16728_ (.A(net349),
    .B(_02371_),
    .X(_02372_));
 inv_2 _16729_ (.A(_02372_),
    .Y(_02373_));
 xnor2_1 _16730_ (.A(_11463_),
    .B(_02357_),
    .Y(_02374_));
 mux2_1 _16731_ (.A0(_02371_),
    .A1(_02373_),
    .S(_11456_),
    .X(_02375_));
 xor2_1 _16732_ (.A(_02362_),
    .B(_02368_),
    .X(_02376_));
 xnor2_1 _16733_ (.A(_02358_),
    .B(_02376_),
    .Y(_02377_));
 xor2_1 _16734_ (.A(_11456_),
    .B(_02372_),
    .X(_02378_));
 xnor2_1 _16735_ (.A(_02285_),
    .B(_02378_),
    .Y(_02379_));
 nor2_1 _16736_ (.A(_02377_),
    .B(_02379_),
    .Y(_02380_));
 nand2_1 _16737_ (.A(_02377_),
    .B(_02379_),
    .Y(_02381_));
 and3b_1 _16738_ (.A_N(_02380_),
    .B(_02381_),
    .C(net468),
    .X(_02382_));
 or4_1 _16739_ (.A(_02339_),
    .B(_02344_),
    .C(_02354_),
    .D(_02382_),
    .X(_02383_));
 mux2_1 _16740_ (.A0(\digitop_pav2.aes128_inst.aes128_regs.state2_r[3] ),
    .A1(_02383_),
    .S(net161),
    .X(_00360_));
 a21o_1 _16741_ (.A1(_11252_),
    .A2(_11290_),
    .B1(net246),
    .X(_02384_));
 nor2_1 _16742_ (.A(_11347_),
    .B(_11494_),
    .Y(_02385_));
 a21o_1 _16743_ (.A1(_11277_),
    .A2(_11320_),
    .B1(_11488_),
    .X(_02386_));
 nor2_1 _16744_ (.A(_11265_),
    .B(_11289_),
    .Y(_02387_));
 a31o_1 _16745_ (.A1(net247),
    .A2(_11292_),
    .A3(_11486_),
    .B1(_11387_),
    .X(_02388_));
 or4_1 _16746_ (.A(net227),
    .B(_11283_),
    .C(_11287_),
    .D(_11365_),
    .X(_02389_));
 or3_2 _16747_ (.A(net246),
    .B(_11291_),
    .C(_11293_),
    .X(_02390_));
 o21ai_1 _16748_ (.A1(net241),
    .A2(_11309_),
    .B1(_02390_),
    .Y(_02391_));
 o311a_1 _16749_ (.A1(net233),
    .A2(_02239_),
    .A3(_02385_),
    .B1(_02386_),
    .C1(net252),
    .X(_02392_));
 a311o_1 _16750_ (.A1(net249),
    .A2(_02388_),
    .A3(_02389_),
    .B1(_02392_),
    .C1(_11357_),
    .X(_02393_));
 o21ai_1 _16751_ (.A1(_02319_),
    .A2(_02387_),
    .B1(net253),
    .Y(_02394_));
 o211a_1 _16752_ (.A1(net253),
    .A2(_02391_),
    .B1(_02394_),
    .C1(net226),
    .X(_02395_));
 o221ai_1 _16753_ (.A1(_11242_),
    .A2(_11264_),
    .B1(_11296_),
    .B2(net247),
    .C1(net249),
    .Y(_02396_));
 o311a_1 _16754_ (.A1(net249),
    .A2(_11263_),
    .A3(_11384_),
    .B1(_02396_),
    .C1(net232),
    .X(_02397_));
 o311a_1 _16755_ (.A1(net281),
    .A2(_02395_),
    .A3(_02397_),
    .B1(_02393_),
    .C1(net286),
    .X(_02398_));
 a31o_1 _16756_ (.A1(net242),
    .A2(_11286_),
    .A3(_11314_),
    .B1(_11344_),
    .X(_02399_));
 o21a_1 _16757_ (.A1(_11261_),
    .A2(_11280_),
    .B1(_11494_),
    .X(_02400_));
 o211a_1 _16758_ (.A1(net233),
    .A2(_02400_),
    .B1(_02399_),
    .C1(net249),
    .X(_02401_));
 or3_2 _16759_ (.A(net232),
    .B(_11319_),
    .C(_11320_),
    .X(_02402_));
 a31o_1 _16760_ (.A1(net245),
    .A2(_11277_),
    .A3(_11347_),
    .B1(_02402_),
    .X(_02403_));
 o221a_1 _16761_ (.A1(net242),
    .A2(_11260_),
    .B1(_11329_),
    .B2(_02170_),
    .C1(net228),
    .X(_02404_));
 and3b_1 _16762_ (.A_N(_02404_),
    .B(net252),
    .C(_02403_),
    .X(_02405_));
 a211o_1 _16763_ (.A1(_11262_),
    .A2(_11320_),
    .B1(_02387_),
    .C1(net249),
    .X(_02406_));
 o311a_1 _16764_ (.A1(net252),
    .A2(_11282_),
    .A3(_11332_),
    .B1(_02406_),
    .C1(net225),
    .X(_02407_));
 o211ai_1 _16765_ (.A1(_11289_),
    .A2(_11329_),
    .B1(_02248_),
    .C1(net252),
    .Y(_02408_));
 a211o_1 _16766_ (.A1(_11281_),
    .A2(_02159_),
    .B1(_02169_),
    .C1(net252),
    .X(_02409_));
 a311o_1 _16767_ (.A1(net233),
    .A2(_02408_),
    .A3(_02409_),
    .B1(_11357_),
    .C1(_02407_),
    .X(_02410_));
 o311a_1 _16768_ (.A1(net280),
    .A2(_02401_),
    .A3(_02405_),
    .B1(_02410_),
    .C1(net283),
    .X(_02411_));
 nor2_2 _16769_ (.A(_02398_),
    .B(_02411_),
    .Y(_02412_));
 and2_2 _16770_ (.A(net472),
    .B(_02412_),
    .X(_02413_));
 nor2_1 _16771_ (.A(net1036),
    .B(_07550_),
    .Y(_02414_));
 a31o_1 _16772_ (.A1(\digitop_pav2.sec_inst.shift_in.s4.q[4] ),
    .A2(net683),
    .A3(net577),
    .B1(_11407_),
    .X(_02415_));
 a31o_1 _16773_ (.A1(\digitop_pav2.sec_inst.shift_in.s6.q[4] ),
    .A2(net598),
    .A3(net594),
    .B1(_02415_),
    .X(_02416_));
 a31o_1 _16774_ (.A1(\digitop_pav2.sec_inst.shift_in.s2.q[4] ),
    .A2(net599),
    .A3(_11417_),
    .B1(_02416_),
    .X(_02417_));
 a221o_1 _16775_ (.A1(\digitop_pav2.sec_inst.shift_in.s12.q[4] ),
    .A2(_11426_),
    .B1(_11428_),
    .B2(\digitop_pav2.sec_inst.shift_in.s10.q[4] ),
    .C1(net576),
    .X(_02418_));
 a21o_1 _16776_ (.A1(\digitop_pav2.sec_inst.shift_in.s8.q[4] ),
    .A2(net574),
    .B1(_11433_),
    .X(_02419_));
 o211a_1 _16777_ (.A1(net1123),
    .A2(net717),
    .B1(net601),
    .C1(_02419_),
    .X(_02420_));
 a32o_1 _16778_ (.A1(_02417_),
    .A2(_02418_),
    .A3(_02420_),
    .B1(net603),
    .B2(_08890_),
    .X(_02421_));
 a22o_1 _16779_ (.A1(net1123),
    .A2(_02414_),
    .B1(_02421_),
    .B2(net534),
    .X(_02422_));
 and2_2 _16780_ (.A(net398),
    .B(_02422_),
    .X(_02423_));
 a221o_1 _16781_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[3] ),
    .A2(net185),
    .B1(net163),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[3] ),
    .C1(net177),
    .X(_02424_));
 a21o_1 _16782_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[3] ),
    .A2(net168),
    .B1(_02424_),
    .X(_02425_));
 o21ai_1 _16783_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[3] ),
    .A2(net175),
    .B1(_02425_),
    .Y(_02426_));
 inv_2 _16784_ (.A(_02426_),
    .Y(_02427_));
 or2_2 _16785_ (.A(net349),
    .B(_02426_),
    .X(_02428_));
 a22o_1 _16786_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[12] ),
    .A2(net168),
    .B1(_11445_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[12] ),
    .X(_02429_));
 a211o_1 _16787_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[12] ),
    .A2(net164),
    .B1(net178),
    .C1(_02429_),
    .X(_02430_));
 o21ai_2 _16788_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[12] ),
    .A2(net175),
    .B1(_02430_),
    .Y(_02431_));
 a22o_1 _16789_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[4] ),
    .A2(net164),
    .B1(_11445_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[4] ),
    .X(_02432_));
 a211o_1 _16790_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[4] ),
    .A2(net168),
    .B1(net178),
    .C1(_02432_),
    .X(_02433_));
 o211ai_4 _16791_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[4] ),
    .A2(net175),
    .B1(_02433_),
    .C1(_11441_),
    .Y(_02434_));
 nor2_2 _16792_ (.A(net349),
    .B(_02431_),
    .Y(_02435_));
 and3_1 _16793_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[12] ),
    .B(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_9.Y ),
    .C(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_9.Y ),
    .X(_02436_));
 a221o_1 _16794_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[12] ),
    .A2(net187),
    .B1(net165),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[12] ),
    .C1(net178),
    .X(_02437_));
 o22a_1 _16795_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[12] ),
    .A2(net173),
    .B1(_02436_),
    .B2(_02437_),
    .X(_02438_));
 nand2_2 _16796_ (.A(_11441_),
    .B(_02438_),
    .Y(_02439_));
 o21ai_1 _16797_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[4] ),
    .B1(net440),
    .Y(_02440_));
 a21oi_1 _16798_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[4] ),
    .B1(_02440_),
    .Y(_02441_));
 or2_1 _16799_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[4] ),
    .X(_02442_));
 nand2_1 _16800_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[4] ),
    .Y(_02443_));
 a31o_1 _16801_ (.A1(net428),
    .A2(_02442_),
    .A3(_02443_),
    .B1(_02441_),
    .X(_02444_));
 xnor2_2 _16802_ (.A(_11462_),
    .B(_02428_),
    .Y(_02445_));
 mux2_1 _16803_ (.A0(_02431_),
    .A1(_02435_),
    .S(_02434_),
    .X(_02446_));
 xnor2_1 _16804_ (.A(_02445_),
    .B(_02446_),
    .Y(_02447_));
 xor2_1 _16805_ (.A(_02378_),
    .B(_02439_),
    .X(_02448_));
 nor2_1 _16806_ (.A(_02447_),
    .B(_02448_),
    .Y(_02449_));
 nand2_1 _16807_ (.A(_02447_),
    .B(_02448_),
    .Y(_02450_));
 and3b_1 _16808_ (.A_N(_02449_),
    .B(_02450_),
    .C(net469),
    .X(_02451_));
 or4_1 _16809_ (.A(_02413_),
    .B(_02423_),
    .C(_02444_),
    .D(_02451_),
    .X(_02452_));
 mux2_1 _16810_ (.A0(\digitop_pav2.aes128_inst.aes128_regs.state2_r[4] ),
    .A1(_02452_),
    .S(net161),
    .X(_00361_));
 a21bo_1 _16811_ (.A1(_11282_),
    .A2(_02160_),
    .B1_N(_02164_),
    .X(_02453_));
 a21oi_1 _16812_ (.A1(net222),
    .A2(_02453_),
    .B1(net286),
    .Y(_02454_));
 a21o_1 _16813_ (.A1(_11277_),
    .A2(_11370_),
    .B1(_11344_),
    .X(_02455_));
 a311o_1 _16814_ (.A1(_11331_),
    .A2(_11339_),
    .A3(_11343_),
    .B1(_11366_),
    .C1(net229),
    .X(_02456_));
 a21o_1 _16815_ (.A1(net238),
    .A2(_11275_),
    .B1(net222),
    .X(_02457_));
 o211a_1 _16816_ (.A1(_02228_),
    .A2(_02457_),
    .B1(_02456_),
    .C1(net284),
    .X(_02458_));
 or4_1 _16817_ (.A(_11261_),
    .B(_11275_),
    .C(_11289_),
    .D(_11313_),
    .X(_02459_));
 nand2_1 _16818_ (.A(_11235_),
    .B(_02459_),
    .Y(_02460_));
 a221o_1 _16819_ (.A1(net239),
    .A2(_11276_),
    .B1(_11295_),
    .B2(_11330_),
    .C1(net224),
    .X(_02461_));
 o2bb2a_1 _16820_ (.A1_N(net200),
    .A2_N(_11311_),
    .B1(_02160_),
    .B2(_11281_),
    .X(_02462_));
 o21ba_1 _16821_ (.A1(net246),
    .A2(_11296_),
    .B1_N(_02246_),
    .X(_02463_));
 or2_1 _16822_ (.A(_11495_),
    .B(_02236_),
    .X(_02464_));
 o221a_1 _16823_ (.A1(_11264_),
    .A2(_11281_),
    .B1(_11313_),
    .B2(_02464_),
    .C1(net232),
    .X(_02465_));
 o21a_1 _16824_ (.A1(_02463_),
    .A2(_02465_),
    .B1(net285),
    .X(_02466_));
 nand2_1 _16825_ (.A(net232),
    .B(_11310_),
    .Y(_02467_));
 o221a_1 _16826_ (.A1(_11309_),
    .A2(_02240_),
    .B1(_02325_),
    .B2(_02467_),
    .C1(net283),
    .X(_02468_));
 nand4_1 _16827_ (.A(net229),
    .B(_11277_),
    .C(_11328_),
    .D(_02152_),
    .Y(_02469_));
 o2bb2a_1 _16828_ (.A1_N(net236),
    .A2_N(_11311_),
    .B1(_11282_),
    .B2(_11265_),
    .X(_02470_));
 o211a_1 _16829_ (.A1(net230),
    .A2(_02470_),
    .B1(_02469_),
    .C1(net282),
    .X(_02471_));
 a221o_1 _16830_ (.A1(net243),
    .A2(_11340_),
    .B1(_11367_),
    .B2(_02163_),
    .C1(net228),
    .X(_02472_));
 o311a_1 _16831_ (.A1(net223),
    .A2(_11320_),
    .A3(_02387_),
    .B1(_02472_),
    .C1(net286),
    .X(_02473_));
 or3_1 _16832_ (.A(net253),
    .B(_02471_),
    .C(_02473_),
    .X(_02474_));
 o311a_1 _16833_ (.A1(net249),
    .A2(_02466_),
    .A3(_02468_),
    .B1(_02474_),
    .C1(net281),
    .X(_02475_));
 a211o_1 _16834_ (.A1(_02454_),
    .A2(_02455_),
    .B1(_02458_),
    .C1(net248),
    .X(_02476_));
 a21o_1 _16835_ (.A1(_02227_),
    .A2(_02460_),
    .B1(net231),
    .X(_02477_));
 or3b_1 _16836_ (.A(_11266_),
    .B(net225),
    .C_N(_11342_),
    .X(_02478_));
 o211a_1 _16837_ (.A1(net229),
    .A2(_02462_),
    .B1(_02461_),
    .C1(net284),
    .X(_02479_));
 a311o_1 _16838_ (.A1(net283),
    .A2(_02477_),
    .A3(_02478_),
    .B1(_02479_),
    .C1(net251),
    .X(_02480_));
 a311oi_2 _16839_ (.A1(_11357_),
    .A2(_02476_),
    .A3(_02480_),
    .B1(_11362_),
    .C1(_02475_),
    .Y(_02481_));
 and2_2 _16840_ (.A(net472),
    .B(net160),
    .X(_02482_));
 o21a_1 _16841_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[13] ),
    .A2(net183),
    .B1(net186),
    .X(_02483_));
 a221o_1 _16842_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[13] ),
    .A2(net168),
    .B1(net164),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[13] ),
    .C1(_02483_),
    .X(_02484_));
 o21ai_1 _16843_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[13] ),
    .A2(net175),
    .B1(_02484_),
    .Y(_02485_));
 or2_2 _16844_ (.A(net349),
    .B(_02485_),
    .X(_02486_));
 inv_2 _16845_ (.A(_02486_),
    .Y(_02487_));
 o21a_1 _16846_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[4] ),
    .A2(net183),
    .B1(net186),
    .X(_02488_));
 a221o_1 _16847_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[4] ),
    .A2(net168),
    .B1(net164),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[4] ),
    .C1(_02488_),
    .X(_02489_));
 o21a_1 _16848_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[4] ),
    .A2(net175),
    .B1(_02489_),
    .X(_02490_));
 nand2_2 _16849_ (.A(_11441_),
    .B(_02490_),
    .Y(_02491_));
 a221o_1 _16850_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[13] ),
    .A2(net186),
    .B1(net163),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[13] ),
    .C1(net177),
    .X(_02492_));
 a21o_1 _16851_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[13] ),
    .A2(net168),
    .B1(_02492_),
    .X(_02493_));
 o21ai_2 _16852_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[13] ),
    .A2(net175),
    .B1(_02493_),
    .Y(_02494_));
 o21a_1 _16853_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[5] ),
    .A2(net183),
    .B1(net186),
    .X(_02495_));
 a221o_1 _16854_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[5] ),
    .A2(net168),
    .B1(net164),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[5] ),
    .C1(_02495_),
    .X(_02496_));
 o21a_1 _16855_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[5] ),
    .A2(net175),
    .B1(_02496_),
    .X(_02497_));
 nand2_2 _16856_ (.A(_11441_),
    .B(_02497_),
    .Y(_02498_));
 or2_2 _16857_ (.A(net349),
    .B(_02494_),
    .X(_02499_));
 inv_2 _16858_ (.A(_02499_),
    .Y(_02500_));
 a221o_1 _16859_ (.A1(\digitop_pav2.sec_inst.shift_in.s12.q[5] ),
    .A2(_11426_),
    .B1(_11428_),
    .B2(\digitop_pav2.sec_inst.shift_in.s10.q[5] ),
    .C1(net576),
    .X(_02501_));
 or2_1 _16860_ (.A(net1120),
    .B(net718),
    .X(_02502_));
 a31o_1 _16861_ (.A1(\digitop_pav2.sec_inst.shift_in.s4.q[5] ),
    .A2(net683),
    .A3(net577),
    .B1(net598),
    .X(_02503_));
 a31o_1 _16862_ (.A1(\digitop_pav2.sec_inst.shift_in.s2.q[5] ),
    .A2(_11397_),
    .A3(net599),
    .B1(_02503_),
    .X(_02504_));
 a21o_1 _16863_ (.A1(\digitop_pav2.sec_inst.shift_in.s6.q[5] ),
    .A2(_11420_),
    .B1(net596),
    .X(_02505_));
 a31o_1 _16864_ (.A1(\digitop_pav2.sec_inst.shift_in.s8.q[5] ),
    .A2(_11404_),
    .A3(net574),
    .B1(_11406_),
    .X(_02506_));
 a31o_1 _16865_ (.A1(net682),
    .A2(_02504_),
    .A3(_02505_),
    .B1(_02506_),
    .X(_02507_));
 a31o_1 _16866_ (.A1(_02501_),
    .A2(_02502_),
    .A3(_02507_),
    .B1(net602),
    .X(_02508_));
 o211a_1 _16867_ (.A1(_08895_),
    .A2(net600),
    .B1(net535),
    .C1(_02508_),
    .X(_02509_));
 o31a_1 _16868_ (.A1(net1036),
    .A2(net1120),
    .A3(net1017),
    .B1(net1255),
    .X(_02510_));
 o21a_2 _16869_ (.A1(_02509_),
    .A2(_02510_),
    .B1(_07519_),
    .X(_02511_));
 o21ai_1 _16870_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[5] ),
    .B1(net440),
    .Y(_02512_));
 a21oi_1 _16871_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[5] ),
    .B1(_02512_),
    .Y(_02513_));
 or2_1 _16872_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[5] ),
    .X(_02514_));
 nand2_1 _16873_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[5] ),
    .Y(_02515_));
 a31o_1 _16874_ (.A1(net428),
    .A2(_02514_),
    .A3(_02515_),
    .B1(_02513_),
    .X(_02516_));
 xnor2_1 _16875_ (.A(_02491_),
    .B(_02498_),
    .Y(_02517_));
 xnor2_1 _16876_ (.A(_02499_),
    .B(_02517_),
    .Y(_02518_));
 xnor2_1 _16877_ (.A(_02439_),
    .B(_02486_),
    .Y(_02519_));
 nor2_1 _16878_ (.A(_02518_),
    .B(_02519_),
    .Y(_02520_));
 nand2_1 _16879_ (.A(_02518_),
    .B(_02519_),
    .Y(_02521_));
 and3b_1 _16880_ (.A_N(_02520_),
    .B(_02521_),
    .C(net469),
    .X(_02522_));
 or4_1 _16881_ (.A(_02482_),
    .B(_02511_),
    .C(_02516_),
    .D(_02522_),
    .X(_02523_));
 mux2_1 _16882_ (.A0(\digitop_pav2.aes128_inst.aes128_regs.state2_r[5] ),
    .A1(_02523_),
    .S(_11204_),
    .X(_00362_));
 nor2_1 _16883_ (.A(_11285_),
    .B(_11329_),
    .Y(_02524_));
 a31o_1 _16884_ (.A1(net241),
    .A2(_11279_),
    .A3(_11308_),
    .B1(_02524_),
    .X(_02525_));
 a21oi_1 _16885_ (.A1(net246),
    .A2(_11282_),
    .B1(_02402_),
    .Y(_02526_));
 a21oi_1 _16886_ (.A1(net231),
    .A2(_02525_),
    .B1(_02526_),
    .Y(_02527_));
 o21ai_1 _16887_ (.A1(_11264_),
    .A2(_11290_),
    .B1(_02390_),
    .Y(_02528_));
 o211a_1 _16888_ (.A1(net238),
    .A2(_02459_),
    .B1(_11376_),
    .C1(net226),
    .X(_02529_));
 a31o_1 _16889_ (.A1(_11262_),
    .A2(_11290_),
    .A3(_11294_),
    .B1(net244),
    .X(_02530_));
 o21ai_1 _16890_ (.A1(_11284_),
    .A2(_11368_),
    .B1(_02530_),
    .Y(_02531_));
 nand2_1 _16891_ (.A(net241),
    .B(_11347_),
    .Y(_02532_));
 nand2_1 _16892_ (.A(net246),
    .B(_11261_),
    .Y(_02533_));
 o211a_1 _16893_ (.A1(_11284_),
    .A2(_11312_),
    .B1(_02533_),
    .C1(net226),
    .X(_02534_));
 a21o_1 _16894_ (.A1(net239),
    .A2(_11276_),
    .B1(_11295_),
    .X(_02535_));
 and3_1 _16895_ (.A(net231),
    .B(_11328_),
    .C(_02384_),
    .X(_02536_));
 a311o_1 _16896_ (.A1(_11279_),
    .A2(_11311_),
    .A3(_11331_),
    .B1(_02165_),
    .C1(net226),
    .X(_02537_));
 a31o_1 _16897_ (.A1(net242),
    .A2(_11278_),
    .A3(_11314_),
    .B1(_02325_),
    .X(_02538_));
 a211o_1 _16898_ (.A1(net231),
    .A2(_02531_),
    .B1(_02529_),
    .C1(net253),
    .X(_02539_));
 o211a_1 _16899_ (.A1(net249),
    .A2(_02527_),
    .B1(_02539_),
    .C1(net281),
    .X(_02540_));
 o211a_1 _16900_ (.A1(net232),
    .A2(_02528_),
    .B1(_02238_),
    .C1(net253),
    .X(_02541_));
 a31o_1 _16901_ (.A1(net231),
    .A2(_02227_),
    .A3(_02532_),
    .B1(_02534_),
    .X(_02542_));
 a211oi_1 _16902_ (.A1(net250),
    .A2(_02542_),
    .B1(_02541_),
    .C1(net281),
    .Y(_02543_));
 a221o_1 _16903_ (.A1(_02176_),
    .A2(_02317_),
    .B1(_02535_),
    .B2(net227),
    .C1(net251),
    .X(_02544_));
 a221o_1 _16904_ (.A1(_11318_),
    .A2(_11484_),
    .B1(_02538_),
    .B2(net227),
    .C1(net248),
    .X(_02545_));
 a21oi_1 _16905_ (.A1(_02544_),
    .A2(_02545_),
    .B1(net280),
    .Y(_02546_));
 a311o_1 _16906_ (.A1(net226),
    .A2(_02255_),
    .A3(_02464_),
    .B1(_02536_),
    .C1(net252),
    .X(_02547_));
 o311a_1 _16907_ (.A1(net231),
    .A2(_02325_),
    .A3(_02524_),
    .B1(_02537_),
    .C1(net252),
    .X(_02548_));
 inv_2 _16908_ (.A(_02548_),
    .Y(_02549_));
 a311o_1 _16909_ (.A1(net281),
    .A2(_02547_),
    .A3(_02549_),
    .B1(_02546_),
    .C1(net285),
    .X(_02550_));
 o311a_2 _16910_ (.A1(net283),
    .A2(_02540_),
    .A3(_02543_),
    .B1(_02550_),
    .C1(_11361_),
    .X(_02551_));
 and2_2 _16911_ (.A(net471),
    .B(_02551_),
    .X(_02552_));
 o22a_1 _16912_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[86] ),
    .A2(_11412_),
    .B1(net596),
    .B2(\digitop_pav2.sec_inst.ld_r.reg96_i[54] ),
    .X(_02553_));
 o211a_1 _16913_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[70] ),
    .A2(_11397_),
    .B1(_11403_),
    .C1(_02553_),
    .X(_02554_));
 a211o_1 _16914_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[38] ),
    .A2(_11404_),
    .B1(_11406_),
    .C1(_02554_),
    .X(_02555_));
 mux2_1 _16915_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[22] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[6] ),
    .S(net598),
    .X(_02556_));
 o221a_1 _16916_ (.A1(net1117),
    .A2(net718),
    .B1(net575),
    .B2(_02556_),
    .C1(net600),
    .X(_02557_));
 a22o_1 _16917_ (.A1(_08900_),
    .A2(net602),
    .B1(_02555_),
    .B2(_02557_),
    .X(_02558_));
 nand2_2 _16918_ (.A(net1255),
    .B(net1017),
    .Y(_02559_));
 o31a_1 _16919_ (.A1(net1036),
    .A2(net1117),
    .A3(net1017),
    .B1(net1259),
    .X(_02560_));
 a21oi_1 _16920_ (.A1(net535),
    .A2(_02558_),
    .B1(_02560_),
    .Y(_02561_));
 nor2_4 _16921_ (.A(_07520_),
    .B(_02561_),
    .Y(_02562_));
 o21ai_1 _16922_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[6] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[6] ),
    .B1(net419),
    .Y(_02563_));
 a21oi_1 _16923_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[6] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[6] ),
    .B1(_02563_),
    .Y(_02564_));
 or2_1 _16924_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[6] ),
    .X(_02565_));
 nand2_1 _16925_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[6] ),
    .Y(_02566_));
 a31o_1 _16926_ (.A1(net433),
    .A2(_02565_),
    .A3(_02566_),
    .B1(_02564_),
    .X(_02567_));
 or3b_1 _16927_ (.A(_02562_),
    .B(_02567_),
    .C_N(net161),
    .X(_02568_));
 o21a_1 _16928_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[5] ),
    .A2(net183),
    .B1(net186),
    .X(_02569_));
 a221o_1 _16929_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[5] ),
    .A2(net168),
    .B1(net164),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[5] ),
    .C1(_02569_),
    .X(_02570_));
 o21a_1 _16930_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[5] ),
    .A2(net175),
    .B1(_02570_),
    .X(_02571_));
 nand2_2 _16931_ (.A(_11441_),
    .B(_02571_),
    .Y(_02572_));
 a22o_1 _16932_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[6] ),
    .A2(net185),
    .B1(net183),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[6] ),
    .X(_02573_));
 a211o_1 _16933_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[6] ),
    .A2(net167),
    .B1(net177),
    .C1(_02573_),
    .X(_02574_));
 o21ai_2 _16934_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[6] ),
    .A2(net175),
    .B1(_02574_),
    .Y(_02575_));
 nor2_2 _16935_ (.A(net348),
    .B(_02575_),
    .Y(_02576_));
 a221o_1 _16936_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[14] ),
    .A2(net184),
    .B1(net166),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[14] ),
    .C1(net176),
    .X(_02577_));
 a21o_1 _16937_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[14] ),
    .A2(net162),
    .B1(_02577_),
    .X(_02578_));
 o21ai_2 _16938_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[14] ),
    .A2(net172),
    .B1(_02578_),
    .Y(_02579_));
 nor2_2 _16939_ (.A(net348),
    .B(_02579_),
    .Y(_02580_));
 a22o_1 _16940_ (.A1(_02576_),
    .A2(_02579_),
    .B1(_02580_),
    .B2(_02575_),
    .X(_02581_));
 xor2_1 _16941_ (.A(_02572_),
    .B(_02581_),
    .X(_02582_));
 o21a_1 _16942_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[14] ),
    .A2(_07110_),
    .B1(net184),
    .X(_02583_));
 a221o_1 _16943_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[14] ),
    .A2(net167),
    .B1(net163),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[14] ),
    .C1(_02583_),
    .X(_02584_));
 o21ai_1 _16944_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[14] ),
    .A2(net174),
    .B1(_02584_),
    .Y(_02585_));
 or2_1 _16945_ (.A(net348),
    .B(_02585_),
    .X(_02586_));
 inv_2 _16946_ (.A(_02586_),
    .Y(_02587_));
 xnor2_1 _16947_ (.A(_02486_),
    .B(_02586_),
    .Y(_02588_));
 o21ai_1 _16948_ (.A1(_02582_),
    .A2(_02588_),
    .B1(net467),
    .Y(_02589_));
 a21oi_2 _16949_ (.A1(_02582_),
    .A2(_02588_),
    .B1(_02589_),
    .Y(_02590_));
 o32a_1 _16950_ (.A1(_02552_),
    .A2(_02568_),
    .A3(_02590_),
    .B1(net161),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[6] ),
    .X(_00363_));
 o211a_1 _16951_ (.A1(_02160_),
    .A2(_02171_),
    .B1(_02172_),
    .C1(net224),
    .X(_02591_));
 a31o_1 _16952_ (.A1(net227),
    .A2(_02164_),
    .A3(_02390_),
    .B1(_02591_),
    .X(_02592_));
 nor2_1 _16953_ (.A(net227),
    .B(_11487_),
    .Y(_02593_));
 o221a_1 _16954_ (.A1(_11276_),
    .A2(_11484_),
    .B1(_02163_),
    .B2(net239),
    .C1(net228),
    .X(_02594_));
 a21o_1 _16955_ (.A1(_02315_),
    .A2(_02593_),
    .B1(net248),
    .X(_02595_));
 o221a_1 _16956_ (.A1(net251),
    .A2(_02592_),
    .B1(_02594_),
    .B2(_02595_),
    .C1(_11357_),
    .X(_02596_));
 a21o_1 _16957_ (.A1(_11339_),
    .A2(_11379_),
    .B1(_02319_),
    .X(_02597_));
 or3_1 _16958_ (.A(net245),
    .B(_11282_),
    .C(_11283_),
    .X(_02598_));
 a221o_1 _16959_ (.A1(net225),
    .A2(_02597_),
    .B1(_02598_),
    .B2(_02327_),
    .C1(net251),
    .X(_02599_));
 a41o_1 _16960_ (.A1(net231),
    .A2(_11281_),
    .A3(_11331_),
    .A4(_02533_),
    .B1(net248),
    .X(_02600_));
 a31o_1 _16961_ (.A1(_11265_),
    .A2(net226),
    .A3(_02384_),
    .B1(_02600_),
    .X(_02601_));
 a31o_1 _16962_ (.A1(net280),
    .A2(_02599_),
    .A3(_02601_),
    .B1(net285),
    .X(_02602_));
 a31o_1 _16963_ (.A1(net246),
    .A2(_11277_),
    .A3(_11290_),
    .B1(_02231_),
    .X(_02603_));
 nand2_1 _16964_ (.A(_11347_),
    .B(_02159_),
    .Y(_02604_));
 a32o_1 _16965_ (.A1(net225),
    .A2(_02603_),
    .A3(_02604_),
    .B1(_11298_),
    .B2(_11312_),
    .X(_02605_));
 a21oi_1 _16966_ (.A1(net245),
    .A2(_11334_),
    .B1(_02402_),
    .Y(_02606_));
 a31o_1 _16967_ (.A1(net227),
    .A2(_11339_),
    .A3(_11496_),
    .B1(net251),
    .X(_02607_));
 o221a_1 _16968_ (.A1(net248),
    .A2(_02605_),
    .B1(_02606_),
    .B2(_02607_),
    .C1(net280),
    .X(_02608_));
 o21a_1 _16969_ (.A1(_11265_),
    .A2(_11348_),
    .B1(_02248_),
    .X(_02609_));
 o22a_1 _16970_ (.A1(_11317_),
    .A2(_02169_),
    .B1(_02609_),
    .B2(net222),
    .X(_02610_));
 and3_1 _16971_ (.A(net229),
    .B(_11341_),
    .C(_02310_),
    .X(_02611_));
 o21ai_1 _16972_ (.A1(_11282_),
    .A2(_11340_),
    .B1(_11492_),
    .Y(_02612_));
 a21o_1 _16973_ (.A1(net222),
    .A2(_02612_),
    .B1(net250),
    .X(_02613_));
 o221a_1 _16974_ (.A1(net253),
    .A2(_02610_),
    .B1(_02611_),
    .B2(_02613_),
    .C1(_11357_),
    .X(_02614_));
 o32a_2 _16975_ (.A1(net283),
    .A2(_02608_),
    .A3(_02614_),
    .B1(_02596_),
    .B2(_02602_),
    .X(_02615_));
 and2_1 _16976_ (.A(net471),
    .B(_02615_),
    .X(_02616_));
 or2_1 _16977_ (.A(\digitop_pav2.sec_inst.ld_r.reg96_i[71] ),
    .B(_11397_),
    .X(_02617_));
 o211a_1 _16978_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[87] ),
    .A2(_11396_),
    .B1(net596),
    .C1(_02617_),
    .X(_02618_));
 a211o_1 _16979_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[55] ),
    .A2(net598),
    .B1(_11432_),
    .C1(_02618_),
    .X(_02619_));
 o211a_1 _16980_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[39] ),
    .A2(_11433_),
    .B1(_02619_),
    .C1(net575),
    .X(_02620_));
 or2_1 _16981_ (.A(\digitop_pav2.sec_inst.ld_r.reg96_i[7] ),
    .B(net595),
    .X(_02621_));
 o211a_1 _16982_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[23] ),
    .A2(net597),
    .B1(_11429_),
    .C1(_02621_),
    .X(_02622_));
 or4b_1 _16983_ (.A(net603),
    .B(_02620_),
    .C(_02622_),
    .D_N(net716),
    .X(_02623_));
 o221a_1 _16984_ (.A1(_08897_),
    .A2(net600),
    .B1(_10419_),
    .B2(net1114),
    .C1(net534),
    .X(_02624_));
 a22o_1 _16985_ (.A1(net1114),
    .A2(_02414_),
    .B1(_02623_),
    .B2(_02624_),
    .X(_02625_));
 and2_2 _16986_ (.A(_07519_),
    .B(_02625_),
    .X(_02626_));
 o21ai_1 _16987_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[7] ),
    .B1(net430),
    .Y(_02627_));
 a21oi_1 _16988_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[7] ),
    .B1(_02627_),
    .Y(_02628_));
 or2_1 _16989_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[7] ),
    .X(_02629_));
 nand2_1 _16990_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[7] ),
    .Y(_02630_));
 a31o_1 _16991_ (.A1(net415),
    .A2(_02629_),
    .A3(_02630_),
    .B1(_02628_),
    .X(_02631_));
 o21a_1 _16992_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[7] ),
    .A2(net183),
    .B1(net184),
    .X(_02632_));
 a221o_1 _16993_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[7] ),
    .A2(net166),
    .B1(net162),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ),
    .C1(_02632_),
    .X(_02633_));
 o21ai_1 _16994_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ),
    .A2(net174),
    .B1(_02633_),
    .Y(_02634_));
 or2_4 _16995_ (.A(net348),
    .B(_02634_),
    .X(_02635_));
 inv_2 _16996_ (.A(_02635_),
    .Y(_02636_));
 a22o_1 _16997_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[15] ),
    .A2(net162),
    .B1(_11445_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[15] ),
    .X(_02637_));
 a211o_1 _16998_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[15] ),
    .A2(net166),
    .B1(net176),
    .C1(_02637_),
    .X(_02638_));
 o21a_1 _16999_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[15] ),
    .A2(net172),
    .B1(_02638_),
    .X(_02639_));
 o21ai_1 _17000_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[15] ),
    .A2(net172),
    .B1(_02638_),
    .Y(_02640_));
 o21a_1 _17001_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[6] ),
    .A2(net183),
    .B1(net185),
    .X(_02641_));
 a22o_1 _17002_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[6] ),
    .A2(net167),
    .B1(net163),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[6] ),
    .X(_02642_));
 o221a_2 _17003_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[6] ),
    .A2(net174),
    .B1(_02641_),
    .B2(_02642_),
    .C1(_11441_),
    .X(_02643_));
 nand2_4 _17004_ (.A(_11441_),
    .B(_02639_),
    .Y(_02644_));
 inv_2 _17005_ (.A(_02644_),
    .Y(_02645_));
 xnor2_1 _17006_ (.A(_11456_),
    .B(_02586_),
    .Y(_02646_));
 xor2_1 _17007_ (.A(_02635_),
    .B(_02643_),
    .X(_02647_));
 xnor2_1 _17008_ (.A(_02644_),
    .B(_02647_),
    .Y(_02648_));
 nor2_1 _17009_ (.A(_02646_),
    .B(_02648_),
    .Y(_02649_));
 nand2_1 _17010_ (.A(_02646_),
    .B(_02648_),
    .Y(_02650_));
 and3b_1 _17011_ (.A_N(_02649_),
    .B(_02650_),
    .C(net467),
    .X(_02651_));
 or4_1 _17012_ (.A(_02616_),
    .B(_02626_),
    .C(_02631_),
    .D(_02651_),
    .X(_02652_));
 mux2_1 _17013_ (.A0(\digitop_pav2.aes128_inst.aes128_regs.state2_r[7] ),
    .A1(_02652_),
    .S(net161),
    .X(_00364_));
 or3b_1 _17014_ (.A(_07090_),
    .B(net818),
    .C_N(_07342_),
    .X(_02653_));
 o211ai_1 _17015_ (.A1(net1045),
    .A2(_07031_),
    .B1(_07381_),
    .C1(_07409_),
    .Y(_02654_));
 mux2_1 _17016_ (.A0(_08056_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[0] ),
    .S(net1043),
    .X(_02655_));
 mux2_1 _17017_ (.A0(_02655_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[1] ),
    .S(net680),
    .X(_00371_));
 mux2_1 _17018_ (.A0(_08058_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[1] ),
    .S(net1043),
    .X(_02656_));
 mux2_1 _17019_ (.A0(_02656_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[2] ),
    .S(net680),
    .X(_00372_));
 mux2_1 _17020_ (.A0(_08077_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[2] ),
    .S(net1043),
    .X(_02657_));
 mux2_1 _17021_ (.A0(_02657_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[3] ),
    .S(net680),
    .X(_00373_));
 mux2_1 _17022_ (.A0(_08080_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[3] ),
    .S(net1043),
    .X(_02658_));
 mux2_1 _17023_ (.A0(_02658_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[4] ),
    .S(net680),
    .X(_00374_));
 mux2_1 _17024_ (.A0(_08052_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[4] ),
    .S(net1043),
    .X(_02659_));
 mux2_1 _17025_ (.A0(_02659_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[5] ),
    .S(net680),
    .X(_00375_));
 mux2_1 _17026_ (.A0(_08082_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[5] ),
    .S(net1043),
    .X(_02660_));
 mux2_1 _17027_ (.A0(_02660_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[6] ),
    .S(net680),
    .X(_00376_));
 mux2_1 _17028_ (.A0(_08054_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[6] ),
    .S(net1043),
    .X(_02661_));
 mux2_1 _17029_ (.A0(_02661_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[7] ),
    .S(net680),
    .X(_00377_));
 mux2_1 _17030_ (.A0(_08069_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[7] ),
    .S(net1043),
    .X(_02662_));
 mux2_1 _17031_ (.A0(_02662_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[8] ),
    .S(net680),
    .X(_00378_));
 mux2_1 _17032_ (.A0(_08061_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[8] ),
    .S(net1044),
    .X(_02663_));
 mux2_1 _17033_ (.A0(_02663_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[9] ),
    .S(net681),
    .X(_00379_));
 mux2_1 _17034_ (.A0(_08074_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[9] ),
    .S(net1043),
    .X(_02664_));
 mux2_1 _17035_ (.A0(_02664_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[10] ),
    .S(net680),
    .X(_00380_));
 mux2_1 _17036_ (.A0(_08065_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[10] ),
    .S(net1044),
    .X(_02665_));
 mux2_1 _17037_ (.A0(_02665_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[11] ),
    .S(net681),
    .X(_00381_));
 mux2_1 _17038_ (.A0(_08068_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[11] ),
    .S(net1044),
    .X(_02666_));
 mux2_1 _17039_ (.A0(_02666_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[12] ),
    .S(net681),
    .X(_00382_));
 mux2_1 _17040_ (.A0(_08073_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[12] ),
    .S(net1044),
    .X(_02667_));
 mux2_1 _17041_ (.A0(_02667_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[13] ),
    .S(net681),
    .X(_00383_));
 mux2_1 _17042_ (.A0(_08085_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[13] ),
    .S(net1045),
    .X(_02668_));
 mux2_1 _17043_ (.A0(_02668_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[14] ),
    .S(net681),
    .X(_00384_));
 mux2_1 _17044_ (.A0(_08051_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[14] ),
    .S(net1045),
    .X(_02669_));
 mux2_1 _17045_ (.A0(_02669_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[15] ),
    .S(net681),
    .X(_00385_));
 nor2_1 _17046_ (.A(net1043),
    .B(_08060_),
    .Y(_02670_));
 mux2_1 _17047_ (.A0(_02670_),
    .A1(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[0] ),
    .S(net680),
    .X(_00386_));
 a31o_1 _17048_ (.A1(\digitop_pav2.access_inst.access_transceiver0.wcnt_stb_valid ),
    .A2(_07022_),
    .A3(_07371_),
    .B1(_10426_),
    .X(_02671_));
 o31a_1 _17049_ (.A1(\digitop_pav2.access_inst.access_check0.wcnt_check_zero ),
    .A2(net1011),
    .A3(_10427_),
    .B1(net1194),
    .X(_02672_));
 nand2_2 _17050_ (.A(_02671_),
    .B(_02672_),
    .Y(_02673_));
 nand2_1 _17051_ (.A(\digitop_pav2.access_inst.access_ctrl0.tx_proc_rd_stb_i ),
    .B(_07053_),
    .Y(_02674_));
 o21a_1 _17052_ (.A1(\digitop_pav2.access_inst.access_ctrl0.tx_proc_rd_stb_i ),
    .A2(_07053_),
    .B1(net1011),
    .X(_02675_));
 xor2_1 _17053_ (.A(net1081),
    .B(_09305_),
    .X(_02676_));
 o2bb2a_1 _17054_ (.A1_N(_02674_),
    .A2_N(_02675_),
    .B1(_02676_),
    .B2(net1011),
    .X(_02677_));
 mux2_1 _17055_ (.A0(net1640),
    .A1(_02677_),
    .S(_10426_),
    .X(_02678_));
 mux2_1 _17056_ (.A0(_02678_),
    .A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[0] ),
    .S(_02673_),
    .X(_00387_));
 o21ai_1 _17057_ (.A1(net1081),
    .A2(_07510_),
    .B1(net912),
    .Y(_02679_));
 xnor2_1 _17058_ (.A(net1080),
    .B(_02679_),
    .Y(_02680_));
 xnor2_1 _17059_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[1] ),
    .B(_02674_),
    .Y(_02681_));
 mux2_1 _17060_ (.A0(_02680_),
    .A1(_02681_),
    .S(net1011),
    .X(_02682_));
 mux2_1 _17061_ (.A0(\digitop_pav2.access_inst.access_check0.wordcnt_i[0] ),
    .A1(_02682_),
    .S(_10426_),
    .X(_02683_));
 mux2_1 _17062_ (.A0(_02683_),
    .A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[1] ),
    .S(_02673_),
    .X(_00388_));
 o22a_1 _17063_ (.A1(net1079),
    .A2(net912),
    .B1(_07533_),
    .B2(_09305_),
    .X(_02684_));
 xor2_1 _17064_ (.A(net1078),
    .B(_02684_),
    .X(_02685_));
 or3_1 _17065_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[1] ),
    .B(\digitop_pav2.access_inst.access_check0.wordcnt_i[2] ),
    .C(_02674_),
    .X(_02686_));
 o21ai_1 _17066_ (.A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[1] ),
    .A2(_02674_),
    .B1(\digitop_pav2.access_inst.access_check0.wordcnt_i[2] ),
    .Y(_02687_));
 a31o_1 _17067_ (.A1(net1011),
    .A2(_02686_),
    .A3(_02687_),
    .B1(_10427_),
    .X(_02688_));
 a21oi_1 _17068_ (.A1(_07344_),
    .A2(_02685_),
    .B1(_02688_),
    .Y(_02689_));
 a21o_1 _17069_ (.A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[1] ),
    .A2(_10427_),
    .B1(_02689_),
    .X(_02690_));
 mux2_1 _17070_ (.A0(_02690_),
    .A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[2] ),
    .S(_02673_),
    .X(_00389_));
 nand2_1 _17071_ (.A(net1075),
    .B(_07536_),
    .Y(_02691_));
 inv_2 _17072_ (.A(_02691_),
    .Y(_02692_));
 o21ai_1 _17073_ (.A1(_07534_),
    .A2(_08032_),
    .B1(_07510_),
    .Y(_02693_));
 a21oi_2 _17074_ (.A1(net1080),
    .A2(net1078),
    .B1(net1076),
    .Y(_02694_));
 a311o_1 _17075_ (.A1(net1079),
    .A2(net1077),
    .A3(net1075),
    .B1(net912),
    .C1(_02694_),
    .X(_02695_));
 a21o_1 _17076_ (.A1(_07537_),
    .A2(_02691_),
    .B1(_09305_),
    .X(_02696_));
 and4_1 _17077_ (.A(_07344_),
    .B(_02693_),
    .C(_02695_),
    .D(_02696_),
    .X(_02697_));
 nand2_1 _17078_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[3] ),
    .B(_02686_),
    .Y(_02698_));
 or2_1 _17079_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[3] ),
    .B(_02686_),
    .X(_02699_));
 a31o_1 _17080_ (.A1(net1011),
    .A2(_02698_),
    .A3(_02699_),
    .B1(_10427_),
    .X(_02700_));
 a2bb2o_1 _17081_ (.A1_N(_02697_),
    .A2_N(_02700_),
    .B1(\digitop_pav2.access_inst.access_check0.wordcnt_i[2] ),
    .B2(_10427_),
    .X(_02701_));
 mux2_1 _17082_ (.A0(_02701_),
    .A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[3] ),
    .S(_02673_),
    .X(_00390_));
 o2bb2a_1 _17083_ (.A1_N(_07510_),
    .A2_N(_08032_),
    .B1(_02694_),
    .B2(_07528_),
    .X(_02702_));
 o21a_1 _17084_ (.A1(_09305_),
    .A2(_02691_),
    .B1(_02702_),
    .X(_02703_));
 xnor2_1 _17085_ (.A(net1074),
    .B(_02703_),
    .Y(_02704_));
 xnor2_1 _17086_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[4] ),
    .B(_02699_),
    .Y(_02705_));
 mux2_1 _17087_ (.A0(_02704_),
    .A1(_02705_),
    .S(net1011),
    .X(_02706_));
 mux2_1 _17088_ (.A0(\digitop_pav2.access_inst.access_check0.wordcnt_i[3] ),
    .A1(_02706_),
    .S(_10426_),
    .X(_02707_));
 mux2_1 _17089_ (.A0(_02707_),
    .A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[4] ),
    .S(_02673_),
    .X(_00391_));
 nand2_1 _17090_ (.A(_07529_),
    .B(_02691_),
    .Y(_02708_));
 or2_1 _17091_ (.A(_07530_),
    .B(_08032_),
    .X(_02709_));
 o21ai_1 _17092_ (.A1(net1074),
    .A2(_08032_),
    .B1(net1073),
    .Y(_02710_));
 nand2_1 _17093_ (.A(_02709_),
    .B(_02710_),
    .Y(_02711_));
 or3_1 _17094_ (.A(\digitop_pav2.access_inst.access_check0.wordcnt_i[4] ),
    .B(\digitop_pav2.access_inst.access_check0.wordcnt_i[5] ),
    .C(_02699_),
    .X(_02712_));
 o21ai_1 _17095_ (.A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[4] ),
    .A2(_02699_),
    .B1(\digitop_pav2.access_inst.access_check0.wordcnt_i[5] ),
    .Y(_02713_));
 o21ai_1 _17096_ (.A1(net1074),
    .A2(_02692_),
    .B1(net1073),
    .Y(_02714_));
 a21oi_1 _17097_ (.A1(_02708_),
    .A2(_02714_),
    .B1(_09305_),
    .Y(_02715_));
 mux2_1 _17098_ (.A0(net1073),
    .A1(_08043_),
    .S(_02694_),
    .X(_02716_));
 a221o_1 _17099_ (.A1(_07510_),
    .A2(_02711_),
    .B1(_02716_),
    .B2(_07527_),
    .C1(_02715_),
    .X(_02717_));
 a31o_1 _17100_ (.A1(_07343_),
    .A2(_02712_),
    .A3(_02713_),
    .B1(_10427_),
    .X(_02718_));
 a21oi_1 _17101_ (.A1(_07344_),
    .A2(_02717_),
    .B1(_02718_),
    .Y(_02719_));
 a21o_1 _17102_ (.A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[4] ),
    .A2(_10427_),
    .B1(_02719_),
    .X(_02720_));
 mux2_1 _17103_ (.A0(_02720_),
    .A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[5] ),
    .S(_02673_),
    .X(_00392_));
 nand2_1 _17104_ (.A(net1072),
    .B(_02708_),
    .Y(_02721_));
 o21a_1 _17105_ (.A1(_07532_),
    .A2(_02692_),
    .B1(_02721_),
    .X(_02722_));
 nand2_1 _17106_ (.A(\digitop_pav2.access_inst.access_check0.wordptr_i[6] ),
    .B(_02709_),
    .Y(_02723_));
 o21a_1 _17107_ (.A1(_07532_),
    .A2(_08032_),
    .B1(_02723_),
    .X(_02724_));
 and3_1 _17108_ (.A(net1072),
    .B(_07529_),
    .C(_02694_),
    .X(_02725_));
 a21oi_1 _17109_ (.A1(_07529_),
    .A2(_02694_),
    .B1(net1072),
    .Y(_02726_));
 or3_1 _17110_ (.A(net912),
    .B(_02725_),
    .C(_02726_),
    .X(_02727_));
 o221a_1 _17111_ (.A1(_09305_),
    .A2(_02722_),
    .B1(_02724_),
    .B2(_07511_),
    .C1(_02727_),
    .X(_02728_));
 a2bb2o_1 _17112_ (.A1_N(_07340_),
    .A2_N(_02699_),
    .B1(_02712_),
    .B2(\digitop_pav2.access_inst.access_check0.wordcnt_i[6] ),
    .X(_02729_));
 mux2_1 _17113_ (.A0(_02728_),
    .A1(_02729_),
    .S(_07343_),
    .X(_02730_));
 mux2_1 _17114_ (.A0(\digitop_pav2.access_inst.access_check0.wordcnt_i[5] ),
    .A1(_02730_),
    .S(_10426_),
    .X(_02731_));
 mux2_1 _17115_ (.A0(_02731_),
    .A1(\digitop_pav2.access_inst.access_check0.wordcnt_i[6] ),
    .S(_02673_),
    .X(_00393_));
 or4bb_4 _17116_ (.A(\digitop_pav2.access_inst.access_ctrl0.rx_par0_i ),
    .B(net1210),
    .C_N(_07400_),
    .D_N(_07401_),
    .X(_02732_));
 or2_1 _17117_ (.A(_07403_),
    .B(_02732_),
    .X(_02733_));
 mux2_1 _17118_ (.A0(net1072),
    .A1(\digitop_pav2.access_inst.access_transceiver0.rx_par_buf[14] ),
    .S(_02733_),
    .X(_00394_));
 mux2_1 _17119_ (.A0(\digitop_pav2.access_inst.access_transceiver0.rx_par_buf[14] ),
    .A1(\digitop_pav2.access_inst.access_transceiver0.rx_par_buf[15] ),
    .S(_02733_),
    .X(_00395_));
 a221oi_2 _17120_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[0] ),
    .A2(_10420_),
    .B1(net394),
    .B2(_07517_),
    .C1(_10740_),
    .Y(_02734_));
 nand2_4 _17121_ (.A(net416),
    .B(_11446_),
    .Y(_02735_));
 and3_4 _17122_ (.A(_11198_),
    .B(net334),
    .C(_02735_),
    .X(_02736_));
 nand3_4 _17123_ (.A(_11198_),
    .B(net334),
    .C(_02735_),
    .Y(_02737_));
 o21ai_1 _17124_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[0] ),
    .B1(net434),
    .Y(_02738_));
 a21oi_1 _17125_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[0] ),
    .B1(_02738_),
    .Y(_02739_));
 xor2_1 _17126_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[0] ),
    .X(_02740_));
 a211o_1 _17127_ (.A1(net419),
    .A2(_02740_),
    .B1(_02739_),
    .C1(_02737_),
    .X(_02741_));
 a22o_1 _17128_ (.A1(_11452_),
    .A2(_02206_),
    .B1(_02207_),
    .B2(_11451_),
    .X(_02742_));
 xnor2_1 _17129_ (.A(_02635_),
    .B(_02742_),
    .Y(_02743_));
 a22o_1 _17130_ (.A1(_11471_),
    .A2(_02640_),
    .B1(_02645_),
    .B2(_11470_),
    .X(_02744_));
 nand2_1 _17131_ (.A(_02743_),
    .B(_02744_),
    .Y(_02745_));
 or2_1 _17132_ (.A(_02743_),
    .B(_02744_),
    .X(_02746_));
 a31o_1 _17133_ (.A1(net467),
    .A2(_02745_),
    .A3(_02746_),
    .B1(_11440_),
    .X(_02747_));
 xnor2_1 _17134_ (.A(_11471_),
    .B(_02644_),
    .Y(_02748_));
 o32a_1 _17135_ (.A1(_11393_),
    .A2(_02741_),
    .A3(_02747_),
    .B1(_02736_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[0] ),
    .X(_00396_));
 xor2_1 _17136_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[1] ),
    .X(_02749_));
 o21ai_1 _17137_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[1] ),
    .B1(net434),
    .Y(_02750_));
 a21oi_1 _17138_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[1] ),
    .B1(_02750_),
    .Y(_02751_));
 a211o_1 _17139_ (.A1(net420),
    .A2(_02749_),
    .B1(_02751_),
    .C1(_02737_),
    .X(_02752_));
 xor2_1 _17140_ (.A(_02212_),
    .B(_02290_),
    .X(_02753_));
 xnor2_4 _17141_ (.A(_11467_),
    .B(_02635_),
    .Y(_02754_));
 xnor2_1 _17142_ (.A(_02753_),
    .B(_02754_),
    .Y(_02755_));
 xnor2_1 _17143_ (.A(_02196_),
    .B(_02748_),
    .Y(_02756_));
 xnor2_1 _17144_ (.A(_02755_),
    .B(_02756_),
    .Y(_02757_));
 a21o_1 _17145_ (.A1(net467),
    .A2(_02757_),
    .B1(_02192_),
    .X(_02758_));
 o32a_1 _17146_ (.A1(_02182_),
    .A2(_02752_),
    .A3(_02758_),
    .B1(_02736_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[1] ),
    .X(_00397_));
 xor2_1 _17147_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[2] ),
    .X(_02759_));
 o21ai_1 _17148_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[2] ),
    .B1(net435),
    .Y(_02760_));
 a21oi_1 _17149_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[2] ),
    .B1(_02760_),
    .Y(_02761_));
 xnor2_1 _17150_ (.A(_02201_),
    .B(_02357_),
    .Y(_02762_));
 xnor2_1 _17151_ (.A(_02284_),
    .B(_02762_),
    .Y(_02763_));
 nand2_1 _17152_ (.A(_02196_),
    .B(_02299_),
    .Y(_02764_));
 o21ai_1 _17153_ (.A1(_02196_),
    .A2(_02298_),
    .B1(_02764_),
    .Y(_02765_));
 a21boi_1 _17154_ (.A1(_02763_),
    .A2(_02765_),
    .B1_N(net466),
    .Y(_02766_));
 o21a_1 _17155_ (.A1(_02763_),
    .A2(_02765_),
    .B1(_02766_),
    .X(_02767_));
 a2111o_1 _17156_ (.A1(net421),
    .A2(_02759_),
    .B1(_02761_),
    .C1(_02280_),
    .D1(_02737_),
    .X(_02768_));
 o32a_1 _17157_ (.A1(_02265_),
    .A2(_02767_),
    .A3(_02768_),
    .B1(_02736_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[2] ),
    .X(_00398_));
 xor2_1 _17158_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[3] ),
    .X(_02769_));
 o21ai_1 _17159_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[3] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[3] ),
    .B1(net436),
    .Y(_02770_));
 a21oi_1 _17160_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[3] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[3] ),
    .B1(_02770_),
    .Y(_02771_));
 a2111o_1 _17161_ (.A1(net419),
    .A2(_02769_),
    .B1(_02771_),
    .C1(_02354_),
    .D1(_02737_),
    .X(_02772_));
 xnor2_1 _17162_ (.A(_02372_),
    .B(_02428_),
    .Y(_02773_));
 a22o_1 _17163_ (.A1(_02295_),
    .A2(_02634_),
    .B1(_02636_),
    .B2(_02294_),
    .X(_02774_));
 xnor2_1 _17164_ (.A(_02773_),
    .B(_02774_),
    .Y(_02775_));
 mux2_2 _17165_ (.A0(_02639_),
    .A1(_02644_),
    .S(_02368_),
    .X(_02776_));
 xor2_1 _17166_ (.A(_02299_),
    .B(_02776_),
    .X(_02777_));
 o21ai_1 _17167_ (.A1(_02775_),
    .A2(_02777_),
    .B1(net467),
    .Y(_02778_));
 a21oi_2 _17168_ (.A1(_02775_),
    .A2(_02777_),
    .B1(_02778_),
    .Y(_02779_));
 o32a_1 _17169_ (.A1(_02339_),
    .A2(_02772_),
    .A3(_02779_),
    .B1(_02736_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[3] ),
    .X(_00399_));
 xor2_1 _17170_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[4] ),
    .X(_02780_));
 o21ai_1 _17171_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[4] ),
    .B1(net436),
    .Y(_02781_));
 a21oi_1 _17172_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[4] ),
    .B1(_02781_),
    .Y(_02782_));
 xnor2_1 _17173_ (.A(_02362_),
    .B(_02636_),
    .Y(_02783_));
 xor2_1 _17174_ (.A(_02439_),
    .B(_02491_),
    .X(_02784_));
 xnor2_1 _17175_ (.A(_02783_),
    .B(_02784_),
    .Y(_02785_));
 xor2_1 _17176_ (.A(_02435_),
    .B(_02776_),
    .X(_02786_));
 a21boi_1 _17177_ (.A1(_02785_),
    .A2(_02786_),
    .B1_N(net469),
    .Y(_02787_));
 o21a_1 _17178_ (.A1(_02785_),
    .A2(_02786_),
    .B1(_02787_),
    .X(_02788_));
 a2111o_1 _17179_ (.A1(net422),
    .A2(_02780_),
    .B1(_02782_),
    .C1(_02423_),
    .D1(_02737_),
    .X(_02789_));
 o32a_1 _17180_ (.A1(_02413_),
    .A2(_02788_),
    .A3(_02789_),
    .B1(_02736_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[4] ),
    .X(_00400_));
 xor2_1 _17181_ (.A(_02434_),
    .B(_02486_),
    .X(_02790_));
 a22o_1 _17182_ (.A1(_02435_),
    .A2(_02494_),
    .B1(_02500_),
    .B2(_02431_),
    .X(_02791_));
 xnor2_1 _17183_ (.A(_02790_),
    .B(_02791_),
    .Y(_02792_));
 a21boi_1 _17184_ (.A1(_02572_),
    .A2(_02792_),
    .B1_N(net469),
    .Y(_02793_));
 o21a_1 _17185_ (.A1(_02572_),
    .A2(_02792_),
    .B1(_02793_),
    .X(_02794_));
 o21ai_1 _17186_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[5] ),
    .B1(net437),
    .Y(_02795_));
 a21oi_1 _17187_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[5] ),
    .B1(_02795_),
    .Y(_02796_));
 or2_1 _17188_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[5] ),
    .X(_02797_));
 nand2_1 _17189_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[5] ),
    .Y(_02798_));
 a31o_1 _17190_ (.A1(net423),
    .A2(_02797_),
    .A3(_02798_),
    .B1(_02796_),
    .X(_02799_));
 or4_1 _17191_ (.A(_02511_),
    .B(_02737_),
    .C(_02794_),
    .D(_02799_),
    .X(_02800_));
 o22a_1 _17192_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[5] ),
    .A2(_02736_),
    .B1(_02800_),
    .B2(_02482_),
    .X(_00401_));
 or2_1 _17193_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[6] ),
    .X(_02801_));
 nand2_1 _17194_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[6] ),
    .Y(_02802_));
 or2_1 _17195_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[6] ),
    .X(_02803_));
 nand2_1 _17196_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[6] ),
    .Y(_02804_));
 a311o_1 _17197_ (.A1(net418),
    .A2(_02801_),
    .A3(_02802_),
    .B1(_02562_),
    .C1(_02737_),
    .X(_02805_));
 a31o_1 _17198_ (.A1(net432),
    .A2(_02803_),
    .A3(_02804_),
    .B1(_02805_),
    .X(_02806_));
 mux2_1 _17199_ (.A0(_02579_),
    .A1(_02580_),
    .S(_02499_),
    .X(_02807_));
 xor2_1 _17200_ (.A(_02498_),
    .B(_02643_),
    .X(_02808_));
 xnor2_1 _17201_ (.A(_02587_),
    .B(_02808_),
    .Y(_02809_));
 o21ai_1 _17202_ (.A1(_02807_),
    .A2(_02809_),
    .B1(net467),
    .Y(_02810_));
 a21oi_2 _17203_ (.A1(_02807_),
    .A2(_02809_),
    .B1(_02810_),
    .Y(_02811_));
 o32a_1 _17204_ (.A1(_02552_),
    .A2(_02806_),
    .A3(_02811_),
    .B1(_02736_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[6] ),
    .X(_00402_));
 xor2_1 _17205_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[7] ),
    .X(_02812_));
 o21ai_1 _17206_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[7] ),
    .B1(net415),
    .Y(_02813_));
 a21oi_1 _17207_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[7] ),
    .B1(_02813_),
    .Y(_02814_));
 a211o_1 _17208_ (.A1(net430),
    .A2(_02812_),
    .B1(_02814_),
    .C1(_02737_),
    .X(_02815_));
 mux2_1 _17209_ (.A0(_02644_),
    .A1(_02639_),
    .S(_02580_),
    .X(_02816_));
 a22o_1 _17210_ (.A1(_11462_),
    .A2(_02575_),
    .B1(_02576_),
    .B2(_11461_),
    .X(_02817_));
 xnor2_1 _17211_ (.A(_11457_),
    .B(_02817_),
    .Y(_02818_));
 nand2_1 _17212_ (.A(_02816_),
    .B(_02818_),
    .Y(_02819_));
 or2_1 _17213_ (.A(_02816_),
    .B(_02818_),
    .X(_02820_));
 a31o_1 _17214_ (.A1(net466),
    .A2(_02819_),
    .A3(_02820_),
    .B1(_02626_),
    .X(_02821_));
 o32a_1 _17215_ (.A1(_02616_),
    .A2(_02815_),
    .A3(_02821_),
    .B1(_02736_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[7] ),
    .X(_00403_));
 o22a_2 _17216_ (.A1(_07516_),
    .A2(net360),
    .B1(net395),
    .B2(_11192_),
    .X(_02822_));
 nand2_4 _17217_ (.A(net468),
    .B(_11444_),
    .Y(_02823_));
 a21oi_4 _17218_ (.A1(net416),
    .A2(_11444_),
    .B1(_11194_),
    .Y(_02824_));
 and3_4 _17219_ (.A(_02822_),
    .B(_02823_),
    .C(_02824_),
    .X(_02825_));
 nand3_4 _17220_ (.A(_02822_),
    .B(_02823_),
    .C(_02824_),
    .Y(_02826_));
 a22o_1 _17221_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[5] ),
    .A2(net362),
    .B1(net396),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[5] ),
    .X(_02827_));
 a22o_1 _17222_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[13] ),
    .A2(net361),
    .B1(net357),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[13] ),
    .X(_02828_));
 a221o_1 _17223_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[13] ),
    .A2(net404),
    .B1(net389),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[13] ),
    .C1(net396),
    .X(_02829_));
 a221o_1 _17224_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[13] ),
    .A2(net365),
    .B1(net391),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[13] ),
    .C1(_02829_),
    .X(_02830_));
 a211o_1 _17225_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[13] ),
    .A2(net355),
    .B1(_02828_),
    .C1(_02830_),
    .X(_02831_));
 or2_1 _17226_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[13] ),
    .B(net394),
    .X(_02832_));
 a32oi_4 _17227_ (.A1(net353),
    .A2(_02831_),
    .A3(_02832_),
    .B1(_02827_),
    .B2(net465),
    .Y(_02833_));
 a32o_1 _17228_ (.A1(net353),
    .A2(_02831_),
    .A3(_02832_),
    .B1(_02827_),
    .B2(net465),
    .X(_02834_));
 a22o_1 _17229_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[3] ),
    .A2(net363),
    .B1(net397),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[3] ),
    .X(_02835_));
 a221o_1 _17230_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[11] ),
    .A2(net404),
    .B1(net357),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[11] ),
    .C1(net395),
    .X(_02836_));
 a22o_1 _17231_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[11] ),
    .A2(net364),
    .B1(net360),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[11] ),
    .X(_02837_));
 a22o_1 _17232_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[11] ),
    .A2(net391),
    .B1(net389),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[11] ),
    .X(_02838_));
 a211o_1 _17233_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[11] ),
    .A2(net355),
    .B1(_02837_),
    .C1(_02838_),
    .X(_02839_));
 o221a_2 _17234_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[11] ),
    .A2(net394),
    .B1(_02836_),
    .B2(_02839_),
    .C1(net353),
    .X(_02840_));
 a21oi_2 _17235_ (.A1(net452),
    .A2(_02835_),
    .B1(_02840_),
    .Y(_02841_));
 a21o_1 _17236_ (.A1(net452),
    .A2(_02835_),
    .B1(_02840_),
    .X(_02842_));
 a22o_1 _17237_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[1] ),
    .A2(net363),
    .B1(net397),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[1] ),
    .X(_02843_));
 o21a_1 _17238_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[9] ),
    .A2(_07106_),
    .B1(net403),
    .X(_02844_));
 a221o_1 _17239_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[9] ),
    .A2(net388),
    .B1(net354),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[9] ),
    .C1(_02844_),
    .X(_02845_));
 a22o_1 _17240_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[9] ),
    .A2(net391),
    .B1(net356),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[9] ),
    .X(_02846_));
 a221o_1 _17241_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[9] ),
    .A2(net364),
    .B1(net360),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[9] ),
    .C1(_02846_),
    .X(_02847_));
 o221a_2 _17242_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[9] ),
    .A2(net392),
    .B1(_02845_),
    .B2(_02847_),
    .C1(net353),
    .X(_02848_));
 a21oi_4 _17243_ (.A1(net452),
    .A2(_02843_),
    .B1(_02848_),
    .Y(_02849_));
 a21o_2 _17244_ (.A1(net452),
    .A2(_02843_),
    .B1(_02848_),
    .X(_02850_));
 a22o_1 _17245_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[2] ),
    .A2(net363),
    .B1(net397),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[2] ),
    .X(_02851_));
 and2_1 _17246_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ),
    .B(net388),
    .X(_02852_));
 a221o_1 _17247_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[10] ),
    .A2(net365),
    .B1(net354),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[10] ),
    .C1(_02852_),
    .X(_02853_));
 a221o_1 _17248_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[10] ),
    .A2(net403),
    .B1(net361),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ),
    .C1(net396),
    .X(_02854_));
 a221o_1 _17249_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[10] ),
    .A2(net390),
    .B1(net356),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[10] ),
    .C1(_02854_),
    .X(_02855_));
 o221a_1 _17250_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[10] ),
    .A2(net392),
    .B1(_02853_),
    .B2(_02855_),
    .C1(net353),
    .X(_02856_));
 a21oi_1 _17251_ (.A1(net451),
    .A2(_02851_),
    .B1(_02856_),
    .Y(_02857_));
 clkinv_4 _17252_ (.A(net207),
    .Y(_02858_));
 nor2_2 _17253_ (.A(net209),
    .B(net207),
    .Y(_02859_));
 nand2_1 _17254_ (.A(net210),
    .B(_02858_),
    .Y(_02860_));
 a22o_1 _17255_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[0] ),
    .A2(net363),
    .B1(net397),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[0] ),
    .X(_02861_));
 a22o_1 _17256_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[8] ),
    .A2(net364),
    .B1(net389),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[8] ),
    .X(_02862_));
 a221o_1 _17257_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[8] ),
    .A2(net404),
    .B1(net357),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[8] ),
    .C1(net395),
    .X(_02863_));
 a221o_1 _17258_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[8] ),
    .A2(net391),
    .B1(net355),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[8] ),
    .C1(_02863_),
    .X(_02864_));
 a211o_1 _17259_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[8] ),
    .A2(net360),
    .B1(_02862_),
    .C1(_02864_),
    .X(_02865_));
 or2_1 _17260_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[8] ),
    .B(net392),
    .X(_02866_));
 a32o_1 _17261_ (.A1(net353),
    .A2(_02865_),
    .A3(_02866_),
    .B1(_02861_),
    .B2(net449),
    .X(_02867_));
 inv_4 _17262_ (.A(net205),
    .Y(_02868_));
 nor2_1 _17263_ (.A(_02849_),
    .B(net206),
    .Y(_02869_));
 nor2_2 _17264_ (.A(net210),
    .B(_02858_),
    .Y(_02870_));
 nand2_2 _17265_ (.A(net209),
    .B(net207),
    .Y(_02871_));
 nor2_2 _17266_ (.A(_02858_),
    .B(net205),
    .Y(_02872_));
 nand2_4 _17267_ (.A(net207),
    .B(_02868_),
    .Y(_02873_));
 nor2_4 _17268_ (.A(net209),
    .B(_02868_),
    .Y(_02874_));
 nor2_1 _17269_ (.A(_02870_),
    .B(_02872_),
    .Y(_02875_));
 nand2_1 _17270_ (.A(_02871_),
    .B(_02873_),
    .Y(_02876_));
 nor2_1 _17271_ (.A(net209),
    .B(net205),
    .Y(_02877_));
 nand2_1 _17272_ (.A(_02849_),
    .B(_02868_),
    .Y(_02878_));
 nor2_1 _17273_ (.A(net210),
    .B(_02868_),
    .Y(_02879_));
 nor2_2 _17274_ (.A(net198),
    .B(_02874_),
    .Y(_02880_));
 or2_2 _17275_ (.A(net198),
    .B(_02874_),
    .X(_02881_));
 nor2_2 _17276_ (.A(_02858_),
    .B(_02881_),
    .Y(_02882_));
 nor2_1 _17277_ (.A(_02859_),
    .B(_02882_),
    .Y(_02883_));
 nor2_1 _17278_ (.A(net214),
    .B(_02883_),
    .Y(_02884_));
 a22o_2 _17279_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[4] ),
    .A2(net362),
    .B1(net397),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[4] ),
    .X(_02885_));
 a22o_1 _17280_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[12] ),
    .A2(net364),
    .B1(net361),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[12] ),
    .X(_02886_));
 a221o_1 _17281_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[12] ),
    .A2(net404),
    .B1(net389),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[12] ),
    .C1(net396),
    .X(_02887_));
 a221o_1 _17282_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[12] ),
    .A2(net391),
    .B1(net355),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[12] ),
    .C1(_02887_),
    .X(_02888_));
 a211o_2 _17283_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[12] ),
    .A2(net357),
    .B1(_02886_),
    .C1(_02888_),
    .X(_02889_));
 or2_2 _17284_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[12] ),
    .B(net394),
    .X(_02890_));
 a32oi_4 _17285_ (.A1(net352),
    .A2(_02889_),
    .A3(_02890_),
    .B1(_02885_),
    .B2(net450),
    .Y(_02891_));
 a32o_1 _17286_ (.A1(net352),
    .A2(_02889_),
    .A3(_02890_),
    .B1(_02885_),
    .B2(net450),
    .X(_02892_));
 nor2_4 _17287_ (.A(_02858_),
    .B(_02868_),
    .Y(_02893_));
 nand2_2 _17288_ (.A(net207),
    .B(net205),
    .Y(_02894_));
 nor2_2 _17289_ (.A(net207),
    .B(net206),
    .Y(_02895_));
 nand2_4 _17290_ (.A(net214),
    .B(_02868_),
    .Y(_02896_));
 nand2_1 _17291_ (.A(net213),
    .B(_02872_),
    .Y(_02897_));
 nor2_4 _17292_ (.A(_02850_),
    .B(_02858_),
    .Y(_02898_));
 nand2_4 _17293_ (.A(net210),
    .B(net208),
    .Y(_02899_));
 nand2_1 _17294_ (.A(net213),
    .B(_02899_),
    .Y(_02900_));
 or2_1 _17295_ (.A(_02868_),
    .B(net194),
    .X(_02901_));
 nand2_1 _17296_ (.A(_02897_),
    .B(_02901_),
    .Y(_02902_));
 or2_1 _17297_ (.A(net264),
    .B(_02902_),
    .X(_02903_));
 nand2_2 _17298_ (.A(net213),
    .B(_02858_),
    .Y(_02904_));
 nand2_2 _17299_ (.A(net219),
    .B(net205),
    .Y(_02905_));
 nand2_1 _17300_ (.A(net219),
    .B(net208),
    .Y(_02906_));
 inv_2 _17301_ (.A(_02906_),
    .Y(_02907_));
 or2_2 _17302_ (.A(net212),
    .B(_02895_),
    .X(_02908_));
 nor2_2 _17303_ (.A(net208),
    .B(_02878_),
    .Y(_02909_));
 inv_2 _17304_ (.A(_02909_),
    .Y(_02910_));
 or2_2 _17305_ (.A(net216),
    .B(_02909_),
    .X(_02911_));
 nand2_2 _17306_ (.A(_02871_),
    .B(_02894_),
    .Y(_02912_));
 o22a_1 _17307_ (.A1(net199),
    .A2(_02904_),
    .B1(_02911_),
    .B2(_02912_),
    .X(_02913_));
 o22a_1 _17308_ (.A1(_02884_),
    .A2(_02903_),
    .B1(_02913_),
    .B2(net272),
    .X(_02914_));
 a22o_1 _17309_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[6] ),
    .A2(net363),
    .B1(net397),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[6] ),
    .X(_02915_));
 a221o_1 _17310_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[14] ),
    .A2(net403),
    .B1(net354),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[14] ),
    .C1(net395),
    .X(_02916_));
 a22o_1 _17311_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[14] ),
    .A2(net364),
    .B1(net388),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[14] ),
    .X(_02917_));
 a221o_1 _17312_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[14] ),
    .A2(net360),
    .B1(net391),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[14] ),
    .C1(_02917_),
    .X(_02918_));
 a211o_1 _17313_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[14] ),
    .A2(net356),
    .B1(_02916_),
    .C1(_02918_),
    .X(_02919_));
 or2_1 _17314_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[14] ),
    .B(net393),
    .X(_02920_));
 a32oi_4 _17315_ (.A1(net352),
    .A2(_02919_),
    .A3(_02920_),
    .B1(_02915_),
    .B2(net450),
    .Y(_02921_));
 a32o_1 _17316_ (.A1(net352),
    .A2(_02919_),
    .A3(_02920_),
    .B1(_02915_),
    .B2(net450),
    .X(_02922_));
 nor2_4 _17317_ (.A(net207),
    .B(_02868_),
    .Y(_02923_));
 nand2_2 _17318_ (.A(_02858_),
    .B(net206),
    .Y(_02924_));
 nor2_1 _17319_ (.A(_02850_),
    .B(_02924_),
    .Y(_02925_));
 nand2_1 _17320_ (.A(net219),
    .B(_02858_),
    .Y(_02926_));
 nand2_1 _17321_ (.A(net217),
    .B(_02873_),
    .Y(_02927_));
 nand2_4 _17322_ (.A(net221),
    .B(_02849_),
    .Y(_02928_));
 nand2_4 _17323_ (.A(net218),
    .B(_02871_),
    .Y(_02929_));
 and3_1 _17324_ (.A(_02905_),
    .B(_02926_),
    .C(_02928_),
    .X(_02930_));
 nor2_1 _17325_ (.A(_02925_),
    .B(_02930_),
    .Y(_02931_));
 inv_2 _17326_ (.A(_02931_),
    .Y(_02932_));
 or2_1 _17327_ (.A(_02881_),
    .B(_02904_),
    .X(_02933_));
 and2_1 _17328_ (.A(net261),
    .B(_02933_),
    .X(_02934_));
 nor2_2 _17329_ (.A(_02872_),
    .B(_02923_),
    .Y(_02935_));
 nand2_1 _17330_ (.A(_02873_),
    .B(_02924_),
    .Y(_02936_));
 o31a_1 _17331_ (.A1(net218),
    .A2(_02874_),
    .A3(_02935_),
    .B1(net267),
    .X(_02937_));
 a221o_1 _17332_ (.A1(_02932_),
    .A2(_02934_),
    .B1(_02937_),
    .B2(_02930_),
    .C1(net275),
    .X(_02938_));
 o211a_1 _17333_ (.A1(net279),
    .A2(_02914_),
    .B1(net203),
    .C1(_02938_),
    .X(_02939_));
 a22o_1 _17334_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[7] ),
    .A2(net363),
    .B1(net397),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[7] ),
    .X(_02940_));
 a22o_1 _17335_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[15] ),
    .A2(net360),
    .B1(net356),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[15] ),
    .X(_02941_));
 a221o_1 _17336_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[15] ),
    .A2(net403),
    .B1(net388),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[15] ),
    .C1(net395),
    .X(_02942_));
 a221o_1 _17337_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[15] ),
    .A2(net364),
    .B1(net391),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[15] ),
    .C1(_02942_),
    .X(_02943_));
 a211o_1 _17338_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[15] ),
    .A2(net354),
    .B1(_02941_),
    .C1(_02943_),
    .X(_02944_));
 or2_1 _17339_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[15] ),
    .B(net393),
    .X(_02945_));
 a32oi_4 _17340_ (.A1(net350),
    .A2(_02944_),
    .A3(_02945_),
    .B1(_02940_),
    .B2(net444),
    .Y(_02946_));
 a32o_1 _17341_ (.A1(net350),
    .A2(_02944_),
    .A3(_02945_),
    .B1(_02940_),
    .B2(net445),
    .X(_02947_));
 and3_1 _17342_ (.A(net219),
    .B(_02860_),
    .C(_02935_),
    .X(_02948_));
 nor2_1 _17343_ (.A(net210),
    .B(net208),
    .Y(_02949_));
 nor2_1 _17344_ (.A(_02896_),
    .B(net197),
    .Y(_02950_));
 o21ai_1 _17345_ (.A1(_02948_),
    .A2(_02950_),
    .B1(net269),
    .Y(_02951_));
 a221o_1 _17346_ (.A1(_02881_),
    .A2(_02907_),
    .B1(net197),
    .B2(net213),
    .C1(net270),
    .X(_02952_));
 a21oi_1 _17347_ (.A1(_02951_),
    .A2(_02952_),
    .B1(net275),
    .Y(_02953_));
 o21ai_1 _17348_ (.A1(net198),
    .A2(_02876_),
    .B1(net214),
    .Y(_02954_));
 nand3_1 _17349_ (.A(net272),
    .B(_02911_),
    .C(_02954_),
    .Y(_02955_));
 o21ai_1 _17350_ (.A1(net220),
    .A2(_02909_),
    .B1(net263),
    .Y(_02956_));
 and2_1 _17351_ (.A(net209),
    .B(_02895_),
    .X(_02957_));
 a211o_1 _17352_ (.A1(_02849_),
    .A2(_02893_),
    .B1(_02956_),
    .C1(_02957_),
    .X(_02958_));
 a31o_1 _17353_ (.A1(net276),
    .A2(_02955_),
    .A3(_02958_),
    .B1(net204),
    .X(_02959_));
 o21ai_1 _17354_ (.A1(_02953_),
    .A2(_02959_),
    .B1(net257),
    .Y(_02960_));
 nor2_1 _17355_ (.A(net207),
    .B(_02880_),
    .Y(_02961_));
 o221a_1 _17356_ (.A1(net219),
    .A2(_02882_),
    .B1(_02929_),
    .B2(_02961_),
    .C1(net262),
    .X(_02962_));
 nand2_4 _17357_ (.A(net214),
    .B(net210),
    .Y(_02963_));
 inv_2 _17358_ (.A(_02963_),
    .Y(_02964_));
 nand2_1 _17359_ (.A(net212),
    .B(_02871_),
    .Y(_02965_));
 nor2_1 _17360_ (.A(net218),
    .B(_02893_),
    .Y(_02966_));
 nand2_2 _17361_ (.A(net211),
    .B(_02894_),
    .Y(_02967_));
 o221a_1 _17362_ (.A1(_02928_),
    .A2(_02936_),
    .B1(_02967_),
    .B2(_02881_),
    .C1(net270),
    .X(_02968_));
 o21a_1 _17363_ (.A1(_02962_),
    .A2(_02968_),
    .B1(net278),
    .X(_02969_));
 or2_1 _17364_ (.A(net219),
    .B(_02925_),
    .X(_02970_));
 inv_2 _17365_ (.A(_02970_),
    .Y(_02971_));
 nand2_1 _17366_ (.A(net210),
    .B(_02872_),
    .Y(_02972_));
 and2_1 _17367_ (.A(_02971_),
    .B(_02972_),
    .X(_02973_));
 inv_2 _17368_ (.A(_02973_),
    .Y(_02974_));
 o21ai_1 _17369_ (.A1(_02879_),
    .A2(_02911_),
    .B1(net272),
    .Y(_02975_));
 or3_1 _17370_ (.A(net212),
    .B(net198),
    .C(_02893_),
    .X(_02976_));
 o31a_1 _17371_ (.A1(net218),
    .A2(_02877_),
    .A3(_02923_),
    .B1(_02976_),
    .X(_02977_));
 o221a_1 _17372_ (.A1(_02973_),
    .A2(_02975_),
    .B1(_02977_),
    .B2(net272),
    .C1(net275),
    .X(_02978_));
 o21a_1 _17373_ (.A1(_02969_),
    .A2(_02978_),
    .B1(_02921_),
    .X(_02979_));
 nand2_2 _17374_ (.A(net218),
    .B(_02899_),
    .Y(_02980_));
 nor2_2 _17375_ (.A(net213),
    .B(net206),
    .Y(_02981_));
 nand2_1 _17376_ (.A(_02899_),
    .B(_02981_),
    .Y(_02982_));
 nand2_1 _17377_ (.A(_02873_),
    .B(_02899_),
    .Y(_02983_));
 nand2_1 _17378_ (.A(net216),
    .B(_02983_),
    .Y(_02984_));
 and2_1 _17379_ (.A(net214),
    .B(_02983_),
    .X(_02985_));
 o221a_1 _17380_ (.A1(net198),
    .A2(_02904_),
    .B1(_02964_),
    .B2(_02873_),
    .C1(net267),
    .X(_02986_));
 a311o_1 _17381_ (.A1(_02934_),
    .A2(_02982_),
    .A3(_02984_),
    .B1(_02986_),
    .C1(_02833_),
    .X(_02987_));
 o21a_1 _17382_ (.A1(_02877_),
    .A2(_02980_),
    .B1(_02937_),
    .X(_02988_));
 or2_1 _17383_ (.A(_02898_),
    .B(net197),
    .X(_02989_));
 nor2_1 _17384_ (.A(_02898_),
    .B(net197),
    .Y(_02990_));
 nor2_1 _17385_ (.A(_02893_),
    .B(_02989_),
    .Y(_02991_));
 inv_2 _17386_ (.A(_02991_),
    .Y(_02992_));
 a311o_1 _17387_ (.A1(net261),
    .A2(_02896_),
    .A3(_02992_),
    .B1(_02988_),
    .C1(net274),
    .X(_02993_));
 a31o_1 _17388_ (.A1(net204),
    .A2(_02987_),
    .A3(_02993_),
    .B1(net256),
    .X(_02994_));
 o221a_4 _17389_ (.A1(_02939_),
    .A2(_02960_),
    .B1(_02979_),
    .B2(_02994_),
    .C1(_11361_),
    .X(_02995_));
 and2_2 _17390_ (.A(net471),
    .B(_02995_),
    .X(_02996_));
 o21ai_1 _17391_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[8] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[8] ),
    .B1(net439),
    .Y(_02997_));
 a21oi_1 _17392_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[8] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[8] ),
    .B1(_02997_),
    .Y(_02998_));
 xor2_1 _17393_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[8] ),
    .X(_02999_));
 a211o_1 _17394_ (.A1(net425),
    .A2(_02999_),
    .B1(_02998_),
    .C1(_02826_),
    .X(_03000_));
 and2_1 _17395_ (.A(net1036),
    .B(_08131_),
    .X(_03001_));
 or2_1 _17396_ (.A(_07550_),
    .B(_03001_),
    .X(_03002_));
 a21o_1 _17397_ (.A1(net1153),
    .A2(_07079_),
    .B1(_03002_),
    .X(_03003_));
 or3_2 _17398_ (.A(\digitop_pav2.sec_inst.shift_in.st[0] ),
    .B(\digitop_pav2.sec_inst.shift_in.st[4] ),
    .C(\digitop_pav2.sec_inst.shift_in.st[1] ),
    .X(_03004_));
 nor2_1 _17399_ (.A(_11400_),
    .B(_03004_),
    .Y(_03005_));
 or2_1 _17400_ (.A(_11400_),
    .B(_03004_),
    .X(_03006_));
 a31o_1 _17401_ (.A1(\digitop_pav2.sec_inst.shift_in.s1.q[0] ),
    .A2(_11417_),
    .A3(net593),
    .B1(_11404_),
    .X(_03007_));
 or3b_4 _17402_ (.A(\digitop_pav2.sec_inst.shift_in.st[0] ),
    .B(\digitop_pav2.sec_inst.shift_in.st[4] ),
    .C_N(\digitop_pav2.sec_inst.shift_in.st[1] ),
    .X(_03008_));
 nor2_1 _17403_ (.A(_11400_),
    .B(_03008_),
    .Y(_03009_));
 or2_1 _17404_ (.A(_11400_),
    .B(_03008_),
    .X(_03010_));
 and3_1 _17405_ (.A(\digitop_pav2.sec_inst.shift_in.s3.q[0] ),
    .B(net683),
    .C(_03010_),
    .X(_03011_));
 nor2_1 _17406_ (.A(_11418_),
    .B(_03004_),
    .Y(_03012_));
 or2_1 _17407_ (.A(_11418_),
    .B(_03004_),
    .X(_03013_));
 a31o_1 _17408_ (.A1(\digitop_pav2.sec_inst.shift_in.s5.q[0] ),
    .A2(net597),
    .A3(net591),
    .B1(_03011_),
    .X(_03014_));
 nor2_4 _17409_ (.A(_11418_),
    .B(_03008_),
    .Y(_03015_));
 o21ai_1 _17410_ (.A1(_11418_),
    .A2(_03008_),
    .B1(\digitop_pav2.sec_inst.shift_in.s7.q[0] ),
    .Y(_03016_));
 a2bb2o_1 _17411_ (.A1_N(_03007_),
    .A2_N(_03014_),
    .B1(_03016_),
    .B2(_11404_),
    .X(_03017_));
 nor2_1 _17412_ (.A(_11423_),
    .B(_03004_),
    .Y(_03018_));
 o21a_1 _17413_ (.A1(_07235_),
    .A2(net590),
    .B1(net595),
    .X(_03019_));
 nor2_1 _17414_ (.A(_11423_),
    .B(_03008_),
    .Y(_03020_));
 or2_4 _17415_ (.A(_11423_),
    .B(_03008_),
    .X(_03021_));
 a21oi_1 _17416_ (.A1(\digitop_pav2.sec_inst.shift_in.s11.q[0] ),
    .A2(_03021_),
    .B1(net595),
    .Y(_03022_));
 o32a_1 _17417_ (.A1(net575),
    .A2(_03019_),
    .A3(_03022_),
    .B1(net716),
    .B2(_07079_),
    .X(_03023_));
 o211ai_1 _17418_ (.A1(_11406_),
    .A2(_03017_),
    .B1(_03023_),
    .C1(net601),
    .Y(_03024_));
 o211ai_2 _17419_ (.A1(_08903_),
    .A2(net600),
    .B1(net535),
    .C1(_03024_),
    .Y(_03025_));
 a21oi_4 _17420_ (.A1(_03003_),
    .A2(_03025_),
    .B1(_07520_),
    .Y(_03026_));
 a22o_1 _17421_ (.A1(_11452_),
    .A2(_11466_),
    .B1(_11467_),
    .B2(_11451_),
    .X(_03027_));
 xnor2_1 _17422_ (.A(_02644_),
    .B(_03027_),
    .Y(_03028_));
 or2_1 _17423_ (.A(_02208_),
    .B(_03028_),
    .X(_03029_));
 nand2_1 _17424_ (.A(_02208_),
    .B(_03028_),
    .Y(_03030_));
 a31o_1 _17425_ (.A1(net468),
    .A2(_03029_),
    .A3(_03030_),
    .B1(_03026_),
    .X(_03031_));
 o32a_1 _17426_ (.A1(_02996_),
    .A2(_03000_),
    .A3(_03031_),
    .B1(_02825_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[8] ),
    .X(_00404_));
 or2_2 _17427_ (.A(net198),
    .B(_02923_),
    .X(_03032_));
 or2_1 _17428_ (.A(net199),
    .B(net194),
    .X(_03033_));
 o21ai_1 _17429_ (.A1(net194),
    .A2(_03032_),
    .B1(net259),
    .Y(_03034_));
 a31oi_1 _17430_ (.A1(_02894_),
    .A2(net194),
    .A3(_02910_),
    .B1(_03034_),
    .Y(_03035_));
 o211a_1 _17431_ (.A1(_02870_),
    .A2(_02935_),
    .B1(_02963_),
    .C1(net265),
    .X(_03036_));
 nor2_1 _17432_ (.A(net207),
    .B(_02881_),
    .Y(_03037_));
 nand2_1 _17433_ (.A(_02858_),
    .B(_02880_),
    .Y(_03038_));
 or2_1 _17434_ (.A(_02983_),
    .B(_03037_),
    .X(_03039_));
 or2_1 _17435_ (.A(net217),
    .B(_03039_),
    .X(_03040_));
 or2_1 _17436_ (.A(_02859_),
    .B(_02895_),
    .X(_03041_));
 nor2_1 _17437_ (.A(_02879_),
    .B(_02926_),
    .Y(_03042_));
 o21ai_1 _17438_ (.A1(_02912_),
    .A2(_03041_),
    .B1(net218),
    .Y(_03043_));
 or3_1 _17439_ (.A(net211),
    .B(_02859_),
    .C(_02935_),
    .X(_03044_));
 a31o_1 _17440_ (.A1(net265),
    .A2(_02933_),
    .A3(_03044_),
    .B1(net273),
    .X(_03045_));
 a31o_1 _17441_ (.A1(net259),
    .A2(_03040_),
    .A3(_03043_),
    .B1(_03045_),
    .X(_03046_));
 and3_1 _17442_ (.A(net211),
    .B(net209),
    .C(_02873_),
    .X(_03047_));
 inv_2 _17443_ (.A(_03047_),
    .Y(_03048_));
 o21a_1 _17444_ (.A1(_03042_),
    .A2(_03047_),
    .B1(net260),
    .X(_03049_));
 a41o_1 _17445_ (.A1(net266),
    .A2(_02908_),
    .A3(_02928_),
    .A4(_03040_),
    .B1(_03049_),
    .X(_03050_));
 nand2_1 _17446_ (.A(_02874_),
    .B(_02926_),
    .Y(_03051_));
 a31o_1 _17447_ (.A1(_02897_),
    .A2(_02982_),
    .A3(_03051_),
    .B1(net260),
    .X(_03052_));
 nand2_1 _17448_ (.A(_02896_),
    .B(net197),
    .Y(_03053_));
 and3_1 _17449_ (.A(net260),
    .B(_02905_),
    .C(_03053_),
    .X(_03054_));
 o21ai_1 _17450_ (.A1(_02896_),
    .A2(_02989_),
    .B1(_03054_),
    .Y(_03055_));
 nor2_1 _17451_ (.A(_02882_),
    .B(_03041_),
    .Y(_03056_));
 nor2_1 _17452_ (.A(net219),
    .B(_03056_),
    .Y(_03057_));
 nor2_1 _17453_ (.A(net214),
    .B(_02899_),
    .Y(_03058_));
 or2_1 _17454_ (.A(_02948_),
    .B(_03058_),
    .X(_03059_));
 nor3_1 _17455_ (.A(net262),
    .B(_03057_),
    .C(_03059_),
    .Y(_03060_));
 nand2_1 _17456_ (.A(net212),
    .B(_02870_),
    .Y(_03061_));
 o211a_1 _17457_ (.A1(net212),
    .A2(_02991_),
    .B1(_03061_),
    .C1(net260),
    .X(_03062_));
 o221a_1 _17458_ (.A1(_02874_),
    .A2(_02929_),
    .B1(_02967_),
    .B2(_02898_),
    .C1(net266),
    .X(_03063_));
 nor2_1 _17459_ (.A(net215),
    .B(_02949_),
    .Y(_03064_));
 nand2_1 _17460_ (.A(net211),
    .B(_02923_),
    .Y(_03065_));
 nand2_1 _17461_ (.A(_02963_),
    .B(_03065_),
    .Y(_03066_));
 inv_2 _17462_ (.A(_03066_),
    .Y(_03067_));
 o211a_1 _17463_ (.A1(_02898_),
    .A2(_02908_),
    .B1(_03067_),
    .C1(net278),
    .X(_03068_));
 nand2_2 _17464_ (.A(net209),
    .B(_02936_),
    .Y(_03069_));
 o221a_1 _17465_ (.A1(net205),
    .A2(_02929_),
    .B1(_03069_),
    .B2(net217),
    .C1(net273),
    .X(_03070_));
 nor2_1 _17466_ (.A(_02874_),
    .B(_02906_),
    .Y(_03071_));
 nor3_1 _17467_ (.A(net259),
    .B(_03042_),
    .C(_03071_),
    .Y(_03072_));
 o21ai_1 _17468_ (.A1(net273),
    .A2(_02900_),
    .B1(_03072_),
    .Y(_03073_));
 o311a_1 _17469_ (.A1(net266),
    .A2(_03068_),
    .A3(_03070_),
    .B1(_03073_),
    .C1(_02921_),
    .X(_03074_));
 o311a_1 _17470_ (.A1(net277),
    .A2(_03035_),
    .A3(_03036_),
    .B1(_03046_),
    .C1(net204),
    .X(_03075_));
 a21o_1 _17471_ (.A1(_03052_),
    .A2(_03055_),
    .B1(_02921_),
    .X(_03076_));
 o311a_1 _17472_ (.A1(net204),
    .A2(_03060_),
    .A3(_03062_),
    .B1(_03076_),
    .C1(net277),
    .X(_03077_));
 a41o_1 _17473_ (.A1(net259),
    .A2(_02897_),
    .A3(_02905_),
    .A4(_03038_),
    .B1(net204),
    .X(_03078_));
 o221a_1 _17474_ (.A1(_02921_),
    .A2(_03050_),
    .B1(_03063_),
    .B2(_03078_),
    .C1(net273),
    .X(_03079_));
 o31a_1 _17475_ (.A1(net258),
    .A2(_03077_),
    .A3(_03079_),
    .B1(_11361_),
    .X(_03080_));
 o31a_2 _17476_ (.A1(net256),
    .A2(_03074_),
    .A3(_03075_),
    .B1(_03080_),
    .X(_03081_));
 and2_2 _17477_ (.A(net471),
    .B(_03081_),
    .X(_03082_));
 o21ai_1 _17478_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[9] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[9] ),
    .B1(net429),
    .Y(_03083_));
 a21oi_1 _17479_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[9] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[9] ),
    .B1(_03083_),
    .Y(_03084_));
 or2_1 _17480_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[9] ),
    .X(_03085_));
 nand2_1 _17481_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[9] ),
    .Y(_03086_));
 a31o_1 _17482_ (.A1(net414),
    .A2(_03085_),
    .A3(_03086_),
    .B1(_03084_),
    .X(_03087_));
 nor2_1 _17483_ (.A(_07050_),
    .B(net1106),
    .Y(_03088_));
 a21o_1 _17484_ (.A1(\digitop_pav2.sec_inst.shift_in.s1.q[1] ),
    .A2(net593),
    .B1(_11416_),
    .X(_03089_));
 a21o_1 _17485_ (.A1(\digitop_pav2.sec_inst.shift_in.s3.q[1] ),
    .A2(net592),
    .B1(_11397_),
    .X(_03090_));
 a21o_1 _17486_ (.A1(\digitop_pav2.sec_inst.shift_in.s5.q[1] ),
    .A2(net591),
    .B1(net595),
    .X(_03091_));
 and4_1 _17487_ (.A(net682),
    .B(_03089_),
    .C(_03090_),
    .D(_03091_),
    .X(_03092_));
 nor2_1 _17488_ (.A(net682),
    .B(_03015_),
    .Y(_03093_));
 a211o_1 _17489_ (.A1(\digitop_pav2.sec_inst.shift_in.s7.q[1] ),
    .A2(_03093_),
    .B1(_03092_),
    .C1(_11406_),
    .X(_03094_));
 nor2_1 _17490_ (.A(net597),
    .B(net590),
    .Y(_03095_));
 and2_1 _17491_ (.A(\digitop_pav2.sec_inst.shift_in.s9.q[1] ),
    .B(_03095_),
    .X(_03096_));
 a31o_1 _17492_ (.A1(\digitop_pav2.sec_inst.shift_in.s11.q[1] ),
    .A2(net597),
    .A3(_03021_),
    .B1(net576),
    .X(_03097_));
 o221a_1 _17493_ (.A1(net1106),
    .A2(net718),
    .B1(_03096_),
    .B2(_03097_),
    .C1(net600),
    .X(_03098_));
 a22o_1 _17494_ (.A1(_08911_),
    .A2(net602),
    .B1(_03094_),
    .B2(_03098_),
    .X(_03099_));
 o2bb2a_1 _17495_ (.A1_N(net534),
    .A2_N(_03099_),
    .B1(_03088_),
    .B2(_03002_),
    .X(_03100_));
 nor2_4 _17496_ (.A(_07520_),
    .B(_03100_),
    .Y(_03101_));
 xnor2_1 _17497_ (.A(_02201_),
    .B(_02212_),
    .Y(_03102_));
 xnor2_1 _17498_ (.A(_02748_),
    .B(_03102_),
    .Y(_03103_));
 xnor2_1 _17499_ (.A(_02219_),
    .B(_02291_),
    .Y(_03104_));
 xnor2_1 _17500_ (.A(_03103_),
    .B(_03104_),
    .Y(_03105_));
 nand2_1 _17501_ (.A(net466),
    .B(_03105_),
    .Y(_03106_));
 or4b_1 _17502_ (.A(_03082_),
    .B(_03087_),
    .C(_03101_),
    .D_N(_03106_),
    .X(_03107_));
 mux2_1 _17503_ (.A0(\digitop_pav2.aes128_inst.aes128_regs.state6_r[9] ),
    .A1(_03107_),
    .S(_02825_),
    .X(_00405_));
 o32a_1 _17504_ (.A1(net221),
    .A2(_02883_),
    .A3(_02895_),
    .B1(_02928_),
    .B2(_02893_),
    .X(_03108_));
 nand2_1 _17505_ (.A(net214),
    .B(_02874_),
    .Y(_03109_));
 and3_1 _17506_ (.A(_02871_),
    .B(net271),
    .C(_03109_),
    .X(_03110_));
 o2bb2a_1 _17507_ (.A1_N(_02926_),
    .A2_N(_03110_),
    .B1(_03108_),
    .B2(net271),
    .X(_03111_));
 a31o_1 _17508_ (.A1(net209),
    .A2(net207),
    .A3(net205),
    .B1(net216),
    .X(_03112_));
 nor2_1 _17509_ (.A(_02898_),
    .B(_02935_),
    .Y(_03113_));
 o221a_1 _17510_ (.A1(_02925_),
    .A2(_03112_),
    .B1(_03113_),
    .B2(net221),
    .C1(net263),
    .X(_03114_));
 or3_1 _17511_ (.A(net221),
    .B(net199),
    .C(net197),
    .X(_03115_));
 a31o_1 _17512_ (.A1(net271),
    .A2(_02932_),
    .A3(_03115_),
    .B1(net256),
    .X(_03116_));
 o221a_1 _17513_ (.A1(net258),
    .A2(_03111_),
    .B1(_03114_),
    .B2(_03116_),
    .C1(net279),
    .X(_03117_));
 o22a_1 _17514_ (.A1(net215),
    .A2(_02883_),
    .B1(_02895_),
    .B2(net194),
    .X(_03118_));
 or2_1 _17515_ (.A(_02882_),
    .B(_02957_),
    .X(_03119_));
 a211o_1 _17516_ (.A1(net215),
    .A2(_03119_),
    .B1(_03064_),
    .C1(net264),
    .X(_03120_));
 o211ai_1 _17517_ (.A1(net272),
    .A2(_03118_),
    .B1(_03120_),
    .C1(net256),
    .Y(_03121_));
 a211o_1 _17518_ (.A1(net220),
    .A2(_02870_),
    .B1(net262),
    .C1(_02981_),
    .X(_03122_));
 nor2_1 _17519_ (.A(_02970_),
    .B(_03119_),
    .Y(_03123_));
 a2111o_1 _17520_ (.A1(_02899_),
    .A2(_02971_),
    .B1(_02981_),
    .C1(_03058_),
    .D1(net269),
    .X(_03124_));
 o21ai_1 _17521_ (.A1(_03122_),
    .A2(_03123_),
    .B1(_03124_),
    .Y(_03125_));
 o211a_1 _17522_ (.A1(net257),
    .A2(_03125_),
    .B1(_03121_),
    .C1(net276),
    .X(_03126_));
 nand2_1 _17523_ (.A(_02924_),
    .B(_03064_),
    .Y(_03127_));
 nand2_1 _17524_ (.A(net205),
    .B(_02989_),
    .Y(_03128_));
 nor2_1 _17525_ (.A(_02905_),
    .B(_02990_),
    .Y(_03129_));
 o211a_1 _17526_ (.A1(_02905_),
    .A2(_02990_),
    .B1(net263),
    .C1(_02901_),
    .X(_03130_));
 o211a_1 _17527_ (.A1(net199),
    .A2(_02970_),
    .B1(_03127_),
    .C1(net269),
    .X(_03131_));
 or3_1 _17528_ (.A(net258),
    .B(_03130_),
    .C(_03131_),
    .X(_03132_));
 nor2_1 _17529_ (.A(_02859_),
    .B(_02876_),
    .Y(_03133_));
 nand2_1 _17530_ (.A(net221),
    .B(_03133_),
    .Y(_03134_));
 o21ai_1 _17531_ (.A1(_02870_),
    .A2(_02935_),
    .B1(_03134_),
    .Y(_03135_));
 or3_1 _17532_ (.A(net210),
    .B(net208),
    .C(_02905_),
    .X(_03136_));
 a31o_1 _17533_ (.A1(net221),
    .A2(_02850_),
    .A3(_02872_),
    .B1(net263),
    .X(_03137_));
 a31oi_1 _17534_ (.A1(net213),
    .A2(_02873_),
    .A3(_03128_),
    .B1(_03137_),
    .Y(_03138_));
 a311o_1 _17535_ (.A1(net263),
    .A2(_03135_),
    .A3(_03136_),
    .B1(_03138_),
    .C1(net256),
    .X(_03139_));
 a21oi_1 _17536_ (.A1(net213),
    .A2(net197),
    .B1(_03137_),
    .Y(_03140_));
 o21a_1 _17537_ (.A1(net210),
    .A2(_02967_),
    .B1(net262),
    .X(_03141_));
 a21o_1 _17538_ (.A1(_02929_),
    .A2(_03141_),
    .B1(_02946_),
    .X(_03142_));
 a31o_1 _17539_ (.A1(net213),
    .A2(_02860_),
    .A3(_02935_),
    .B1(net262),
    .X(_03143_));
 a21o_1 _17540_ (.A1(net213),
    .A2(_02898_),
    .B1(_03143_),
    .X(_03144_));
 a31o_1 _17541_ (.A1(net209),
    .A2(_02873_),
    .A3(_02924_),
    .B1(net214),
    .X(_03145_));
 a2bb2o_1 _17542_ (.A1_N(_02884_),
    .A2_N(_03144_),
    .B1(_03145_),
    .B2(_03141_),
    .X(_03146_));
 o221a_1 _17543_ (.A1(_03140_),
    .A2(_03142_),
    .B1(_03146_),
    .B2(net257),
    .C1(net278),
    .X(_03147_));
 a31o_1 _17544_ (.A1(net275),
    .A2(_03132_),
    .A3(_03139_),
    .B1(net204),
    .X(_03148_));
 o32a_4 _17545_ (.A1(_02921_),
    .A2(_03117_),
    .A3(_03126_),
    .B1(_03147_),
    .B2(_03148_),
    .X(_03149_));
 and2_2 _17546_ (.A(net471),
    .B(_03149_),
    .X(_03150_));
 a211o_1 _17547_ (.A1(net1153),
    .A2(net1102),
    .B1(net1017),
    .C1(_03001_),
    .X(_03151_));
 a21o_1 _17548_ (.A1(\digitop_pav2.sec_inst.shift_in.s1.q[2] ),
    .A2(net593),
    .B1(_11416_),
    .X(_03152_));
 a21o_1 _17549_ (.A1(\digitop_pav2.sec_inst.shift_in.s3.q[2] ),
    .A2(net592),
    .B1(_11397_),
    .X(_03153_));
 a21o_1 _17550_ (.A1(\digitop_pav2.sec_inst.shift_in.s5.q[2] ),
    .A2(net591),
    .B1(net595),
    .X(_03154_));
 and4_1 _17551_ (.A(net682),
    .B(_03152_),
    .C(_03153_),
    .D(_03154_),
    .X(_03155_));
 a211o_1 _17552_ (.A1(\digitop_pav2.sec_inst.shift_in.s7.q[2] ),
    .A2(_03093_),
    .B1(_03155_),
    .C1(_11406_),
    .X(_03156_));
 and2_1 _17553_ (.A(\digitop_pav2.sec_inst.shift_in.s9.q[2] ),
    .B(_03095_),
    .X(_03157_));
 a31o_1 _17554_ (.A1(\digitop_pav2.sec_inst.shift_in.s11.q[2] ),
    .A2(net597),
    .A3(_03021_),
    .B1(net576),
    .X(_03158_));
 o221a_1 _17555_ (.A1(net1102),
    .A2(net718),
    .B1(_03157_),
    .B2(_03158_),
    .C1(net600),
    .X(_03159_));
 a22o_1 _17556_ (.A1(_08908_),
    .A2(net602),
    .B1(_03156_),
    .B2(_03159_),
    .X(_03160_));
 a22o_1 _17557_ (.A1(net1255),
    .A2(_03151_),
    .B1(_03160_),
    .B2(net534),
    .X(_03161_));
 and2_2 _17558_ (.A(net398),
    .B(_03161_),
    .X(_03162_));
 o21ai_1 _17559_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[10] ),
    .B1(net431),
    .Y(_03163_));
 a21oi_1 _17560_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[10] ),
    .B1(_03163_),
    .Y(_03164_));
 xor2_1 _17561_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[10] ),
    .X(_03165_));
 a2111o_1 _17562_ (.A1(net416),
    .A2(_03165_),
    .B1(_03164_),
    .C1(_03162_),
    .D1(_02826_),
    .X(_03166_));
 a22o_1 _17563_ (.A1(_02197_),
    .A2(_02294_),
    .B1(_02295_),
    .B2(_02195_),
    .X(_03167_));
 mux2_1 _17564_ (.A0(_02289_),
    .A1(_02291_),
    .S(_02357_),
    .X(_03168_));
 xnor2_1 _17565_ (.A(_02284_),
    .B(_03167_),
    .Y(_03169_));
 o21ai_1 _17566_ (.A1(_03168_),
    .A2(_03169_),
    .B1(net466),
    .Y(_03170_));
 a21oi_2 _17567_ (.A1(_03168_),
    .A2(_03169_),
    .B1(_03170_),
    .Y(_03171_));
 o32a_1 _17568_ (.A1(_03150_),
    .A2(_03166_),
    .A3(_03171_),
    .B1(_02825_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ),
    .X(_00406_));
 o221a_1 _17569_ (.A1(net217),
    .A2(_02882_),
    .B1(_02898_),
    .B2(_02908_),
    .C1(net259),
    .X(_03172_));
 a2bb2o_1 _17570_ (.A1_N(_02961_),
    .A2_N(_02965_),
    .B1(_03032_),
    .B2(net217),
    .X(_03173_));
 a211o_1 _17571_ (.A1(net265),
    .A2(_03173_),
    .B1(_03172_),
    .C1(net273),
    .X(_03174_));
 or2_1 _17572_ (.A(_02935_),
    .B(net197),
    .X(_03175_));
 mux2_1 _17573_ (.A0(_02936_),
    .A1(_03175_),
    .S(_02963_),
    .X(_03176_));
 nor2_1 _17574_ (.A(net265),
    .B(_03176_),
    .Y(_03177_));
 o211a_1 _17575_ (.A1(_02980_),
    .A2(_03032_),
    .B1(_03069_),
    .C1(net265),
    .X(_03178_));
 o311a_1 _17576_ (.A1(net277),
    .A2(_03177_),
    .A3(_03178_),
    .B1(net256),
    .C1(_03174_),
    .X(_03179_));
 o21ai_1 _17577_ (.A1(net213),
    .A2(_02878_),
    .B1(_03044_),
    .Y(_03180_));
 or4b_1 _17578_ (.A(net262),
    .B(_02985_),
    .C(_03180_),
    .D_N(_03065_),
    .X(_03181_));
 a211o_1 _17579_ (.A1(_02878_),
    .A2(_02966_),
    .B1(_03133_),
    .C1(net271),
    .X(_03182_));
 nor2_1 _17580_ (.A(net211),
    .B(_03037_),
    .Y(_03183_));
 o221a_1 _17581_ (.A1(_02971_),
    .A2(_03122_),
    .B1(_03183_),
    .B2(_02956_),
    .C1(net275),
    .X(_03184_));
 a31o_1 _17582_ (.A1(net278),
    .A2(_03181_),
    .A3(_03182_),
    .B1(_03184_),
    .X(_03185_));
 a211o_1 _17583_ (.A1(net258),
    .A2(_03185_),
    .B1(_03179_),
    .C1(net203),
    .X(_03186_));
 o21a_1 _17584_ (.A1(net211),
    .A2(_02961_),
    .B1(_03048_),
    .X(_03187_));
 o21a_1 _17585_ (.A1(_03071_),
    .A2(_03187_),
    .B1(net259),
    .X(_03188_));
 a31o_1 _17586_ (.A1(net265),
    .A2(_02904_),
    .A3(_03032_),
    .B1(_03188_),
    .X(_03189_));
 nand2_1 _17587_ (.A(net277),
    .B(_03189_),
    .Y(_03190_));
 o221a_1 _17588_ (.A1(_02880_),
    .A2(_02929_),
    .B1(_02967_),
    .B2(net198),
    .C1(net259),
    .X(_03191_));
 o221a_1 _17589_ (.A1(_02881_),
    .A2(_02908_),
    .B1(_03175_),
    .B2(net194),
    .C1(net265),
    .X(_03192_));
 o311a_1 _17590_ (.A1(net277),
    .A2(_03191_),
    .A3(_03192_),
    .B1(net256),
    .C1(_03190_),
    .X(_03193_));
 nand2_1 _17591_ (.A(net217),
    .B(_03039_),
    .Y(_03194_));
 or2_1 _17592_ (.A(_02872_),
    .B(_02970_),
    .X(_03195_));
 o221a_1 _17593_ (.A1(_02874_),
    .A2(_02929_),
    .B1(net197),
    .B2(_02896_),
    .C1(net266),
    .X(_03196_));
 a311o_1 _17594_ (.A1(net260),
    .A2(_03194_),
    .A3(_03195_),
    .B1(_03196_),
    .C1(net277),
    .X(_03197_));
 o32a_1 _17595_ (.A1(net269),
    .A2(_02981_),
    .A3(_03058_),
    .B1(_03129_),
    .B2(_02903_),
    .X(_03198_));
 nand2_1 _17596_ (.A(net278),
    .B(_03198_),
    .Y(_03199_));
 a31o_1 _17597_ (.A1(net258),
    .A2(_03197_),
    .A3(_03199_),
    .B1(_03193_),
    .X(_03200_));
 a21bo_2 _17598_ (.A1(net203),
    .A2(_03200_),
    .B1_N(_03186_),
    .X(_03201_));
 and2_2 _17599_ (.A(net473),
    .B(_03201_),
    .X(_03202_));
 o21ai_1 _17600_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[11] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[11] ),
    .B1(net438),
    .Y(_03203_));
 a21oi_1 _17601_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[11] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[11] ),
    .B1(_03203_),
    .Y(_03204_));
 xor2_1 _17602_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[11] ),
    .X(_03205_));
 a21o_1 _17603_ (.A1(\digitop_pav2.sec_inst.shift_in.s5.q[3] ),
    .A2(net591),
    .B1(net595),
    .X(_03206_));
 a21o_1 _17604_ (.A1(\digitop_pav2.sec_inst.shift_in.s3.q[3] ),
    .A2(net592),
    .B1(_11397_),
    .X(_03207_));
 a21o_1 _17605_ (.A1(\digitop_pav2.sec_inst.shift_in.s1.q[3] ),
    .A2(net593),
    .B1(_11416_),
    .X(_03208_));
 nor2_1 _17606_ (.A(net595),
    .B(_03020_),
    .Y(_03209_));
 a221o_1 _17607_ (.A1(\digitop_pav2.sec_inst.shift_in.s9.q[3] ),
    .A2(_03095_),
    .B1(_03209_),
    .B2(\digitop_pav2.sec_inst.shift_in.s11.q[3] ),
    .C1(net575),
    .X(_03210_));
 and3_1 _17608_ (.A(net682),
    .B(_03206_),
    .C(_03208_),
    .X(_03211_));
 a221o_1 _17609_ (.A1(\digitop_pav2.sec_inst.shift_in.s7.q[3] ),
    .A2(_03093_),
    .B1(_03207_),
    .B2(_03211_),
    .C1(_11406_),
    .X(_03212_));
 o211a_1 _17610_ (.A1(net1098),
    .A2(net718),
    .B1(_03210_),
    .C1(_03212_),
    .X(_03213_));
 mux2_1 _17611_ (.A0(_08913_),
    .A1(_03213_),
    .S(net600),
    .X(_03214_));
 nor3_1 _17612_ (.A(net1153),
    .B(_07550_),
    .C(_08118_),
    .Y(_03215_));
 a221o_1 _17613_ (.A1(net1098),
    .A2(_02414_),
    .B1(_03214_),
    .B2(net534),
    .C1(_03215_),
    .X(_03216_));
 and2_2 _17614_ (.A(net398),
    .B(_03216_),
    .X(_03217_));
 xor2_1 _17615_ (.A(_02372_),
    .B(_02644_),
    .X(_03218_));
 mux2_1 _17616_ (.A0(_02361_),
    .A1(_02363_),
    .S(_02299_),
    .X(_03219_));
 xnor2_1 _17617_ (.A(_03218_),
    .B(_03219_),
    .Y(_03220_));
 xnor2_1 _17618_ (.A(_02374_),
    .B(_02428_),
    .Y(_03221_));
 a21boi_1 _17619_ (.A1(_03220_),
    .A2(_03221_),
    .B1_N(net468),
    .Y(_03222_));
 o21a_2 _17620_ (.A1(_03220_),
    .A2(_03221_),
    .B1(_03222_),
    .X(_03223_));
 a2111o_1 _17621_ (.A1(net425),
    .A2(_03205_),
    .B1(_03217_),
    .C1(_02826_),
    .D1(_03204_),
    .X(_03224_));
 o32a_1 _17622_ (.A1(_03202_),
    .A2(_03223_),
    .A3(_03224_),
    .B1(_02825_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[11] ),
    .X(_00407_));
 nor2_1 _17623_ (.A(net221),
    .B(_03133_),
    .Y(_03225_));
 or3_1 _17624_ (.A(_02859_),
    .B(net268),
    .C(_02923_),
    .X(_03226_));
 a21bo_1 _17625_ (.A1(_02879_),
    .A2(net271),
    .B1_N(_03226_),
    .X(_03227_));
 and3_1 _17626_ (.A(_02878_),
    .B(net271),
    .C(_02985_),
    .X(_03228_));
 a221o_1 _17627_ (.A1(net263),
    .A2(_03225_),
    .B1(_03227_),
    .B2(net221),
    .C1(_03228_),
    .X(_03229_));
 o32a_1 _17628_ (.A1(net218),
    .A2(_02877_),
    .A3(_02923_),
    .B1(_02912_),
    .B2(_02911_),
    .X(_03230_));
 nand2_1 _17629_ (.A(net271),
    .B(_03230_),
    .Y(_03231_));
 a211o_1 _17630_ (.A1(net219),
    .A2(net199),
    .B1(net272),
    .C1(_03058_),
    .X(_03232_));
 o211a_1 _17631_ (.A1(_02902_),
    .A2(_03232_),
    .B1(_03231_),
    .C1(net279),
    .X(_03233_));
 a211oi_1 _17632_ (.A1(net275),
    .A2(_03229_),
    .B1(_03233_),
    .C1(net257),
    .Y(_03234_));
 o211a_1 _17633_ (.A1(net214),
    .A2(_03056_),
    .B1(_02954_),
    .C1(net271),
    .X(_03235_));
 or4_1 _17634_ (.A(_02880_),
    .B(net271),
    .C(_02895_),
    .D(_02931_),
    .X(_03236_));
 or3b_1 _17635_ (.A(net279),
    .B(_03235_),
    .C_N(_03236_),
    .X(_03237_));
 a211oi_1 _17636_ (.A1(_02924_),
    .A2(_02964_),
    .B1(_03059_),
    .C1(net263),
    .Y(_03238_));
 o311a_1 _17637_ (.A1(net220),
    .A2(_02879_),
    .A3(_02990_),
    .B1(_03145_),
    .C1(net264),
    .X(_03239_));
 o311a_1 _17638_ (.A1(net276),
    .A2(_03238_),
    .A3(_03239_),
    .B1(net256),
    .C1(_03237_),
    .X(_03240_));
 o21a_1 _17639_ (.A1(net214),
    .A2(_03119_),
    .B1(_02937_),
    .X(_03241_));
 a31o_1 _17640_ (.A1(_02896_),
    .A2(_02912_),
    .A3(_02963_),
    .B1(net272),
    .X(_03242_));
 or3b_1 _17641_ (.A(net279),
    .B(_03241_),
    .C_N(_03242_),
    .X(_03243_));
 o211a_1 _17642_ (.A1(_02895_),
    .A2(_03112_),
    .B1(_02904_),
    .C1(net272),
    .X(_03244_));
 or2_1 _17643_ (.A(_02898_),
    .B(_03127_),
    .X(_03245_));
 or2_1 _17644_ (.A(net270),
    .B(_03066_),
    .X(_03246_));
 a311o_1 _17645_ (.A1(net263),
    .A2(_03067_),
    .A3(_03245_),
    .B1(_03244_),
    .C1(net276),
    .X(_03247_));
 o221a_1 _17646_ (.A1(net194),
    .A2(_02923_),
    .B1(_02929_),
    .B2(net205),
    .C1(net267),
    .X(_03248_));
 a311o_1 _17647_ (.A1(_02875_),
    .A2(net261),
    .A3(_02911_),
    .B1(_03248_),
    .C1(net277),
    .X(_03249_));
 o221a_1 _17648_ (.A1(_02898_),
    .A2(_02908_),
    .B1(_02965_),
    .B2(_02874_),
    .C1(net267),
    .X(_03250_));
 o221a_1 _17649_ (.A1(_02893_),
    .A2(_02963_),
    .B1(_02980_),
    .B2(net198),
    .C1(net261),
    .X(_03251_));
 o311a_1 _17650_ (.A1(net274),
    .A2(_03250_),
    .A3(_03251_),
    .B1(net256),
    .C1(_03249_),
    .X(_03252_));
 a311o_1 _17651_ (.A1(net258),
    .A2(_03243_),
    .A3(_03247_),
    .B1(_03252_),
    .C1(_02921_),
    .X(_03253_));
 o31a_4 _17652_ (.A1(net203),
    .A2(_03234_),
    .A3(_03240_),
    .B1(_03253_),
    .X(_03254_));
 and2_2 _17653_ (.A(net473),
    .B(_03254_),
    .X(_03255_));
 o21ai_1 _17654_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[12] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[12] ),
    .B1(net438),
    .Y(_03256_));
 a21oi_1 _17655_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[12] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[12] ),
    .B1(_03256_),
    .Y(_03257_));
 xor2_1 _17656_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[12] ),
    .X(_03258_));
 a21oi_1 _17657_ (.A1(net1153),
    .A2(net1035),
    .B1(_03002_),
    .Y(_03259_));
 a21o_1 _17658_ (.A1(\digitop_pav2.sec_inst.shift_in.s5.q[4] ),
    .A2(net591),
    .B1(net595),
    .X(_03260_));
 a21o_1 _17659_ (.A1(\digitop_pav2.sec_inst.shift_in.s3.q[4] ),
    .A2(net592),
    .B1(_11397_),
    .X(_03261_));
 a21o_1 _17660_ (.A1(\digitop_pav2.sec_inst.shift_in.s1.q[4] ),
    .A2(_03006_),
    .B1(_11416_),
    .X(_03262_));
 a221o_1 _17661_ (.A1(\digitop_pav2.sec_inst.shift_in.s9.q[4] ),
    .A2(_03095_),
    .B1(_03209_),
    .B2(\digitop_pav2.sec_inst.shift_in.s11.q[4] ),
    .C1(net575),
    .X(_03263_));
 or2_1 _17662_ (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[12] ),
    .B(net718),
    .X(_03264_));
 and3_1 _17663_ (.A(net682),
    .B(_03260_),
    .C(_03262_),
    .X(_03265_));
 a221o_1 _17664_ (.A1(\digitop_pav2.sec_inst.shift_in.s7.q[4] ),
    .A2(_03093_),
    .B1(_03261_),
    .B2(_03265_),
    .C1(_11406_),
    .X(_03266_));
 a31o_1 _17665_ (.A1(_03263_),
    .A2(_03264_),
    .A3(_03266_),
    .B1(net602),
    .X(_03267_));
 o211a_1 _17666_ (.A1(_08909_),
    .A2(net600),
    .B1(net534),
    .C1(_03267_),
    .X(_03268_));
 o21a_4 _17667_ (.A1(_03259_),
    .A2(_03268_),
    .B1(net398),
    .X(_03269_));
 mux2_1 _17668_ (.A0(_02438_),
    .A1(_02439_),
    .S(_02434_),
    .X(_03270_));
 xnor2_1 _17669_ (.A(_02776_),
    .B(_03270_),
    .Y(_03271_));
 xor2_1 _17670_ (.A(_02445_),
    .B(_02491_),
    .X(_03272_));
 a21boi_1 _17671_ (.A1(_03271_),
    .A2(_03272_),
    .B1_N(net469),
    .Y(_03273_));
 o21a_2 _17672_ (.A1(_03271_),
    .A2(_03272_),
    .B1(_03273_),
    .X(_03274_));
 a2111o_1 _17673_ (.A1(net425),
    .A2(_03258_),
    .B1(_03269_),
    .C1(_02826_),
    .D1(_03257_),
    .X(_03275_));
 o32a_1 _17674_ (.A1(_03255_),
    .A2(_03274_),
    .A3(_03275_),
    .B1(_02825_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[12] ),
    .X(_00408_));
 o211a_1 _17675_ (.A1(net198),
    .A2(_02980_),
    .B1(_02963_),
    .C1(net267),
    .X(_03276_));
 a21bo_1 _17676_ (.A1(_02926_),
    .A2(_03128_),
    .B1_N(_03136_),
    .X(_03277_));
 o311a_1 _17677_ (.A1(net218),
    .A2(_02912_),
    .A3(_03037_),
    .B1(_03112_),
    .C1(net267),
    .X(_03278_));
 o22a_1 _17678_ (.A1(_02893_),
    .A2(_02928_),
    .B1(_02984_),
    .B2(_02877_),
    .X(_03279_));
 nor2_1 _17679_ (.A(net267),
    .B(_03279_),
    .Y(_03280_));
 a211o_1 _17680_ (.A1(net261),
    .A2(_03277_),
    .B1(_03276_),
    .C1(net277),
    .X(_03281_));
 o311a_1 _17681_ (.A1(net274),
    .A2(_03278_),
    .A3(_03280_),
    .B1(_03281_),
    .C1(_02921_),
    .X(_03282_));
 o22a_1 _17682_ (.A1(net211),
    .A2(net198),
    .B1(_02896_),
    .B2(_02898_),
    .X(_03283_));
 a211o_1 _17683_ (.A1(_02928_),
    .A2(_03048_),
    .B1(net260),
    .C1(_02923_),
    .X(_03284_));
 o311a_1 _17684_ (.A1(net266),
    .A2(_03071_),
    .A3(_03283_),
    .B1(_03284_),
    .C1(net273),
    .X(_03285_));
 inv_2 _17685_ (.A(_03285_),
    .Y(_03286_));
 a21oi_1 _17686_ (.A1(_02899_),
    .A2(_02966_),
    .B1(_03226_),
    .Y(_03287_));
 a311o_1 _17687_ (.A1(net268),
    .A2(_03038_),
    .A3(_03195_),
    .B1(_03287_),
    .C1(net273),
    .X(_03288_));
 a311o_1 _17688_ (.A1(net204),
    .A2(_03286_),
    .A3(_03288_),
    .B1(net258),
    .C1(_03282_),
    .X(_03289_));
 o21a_1 _17689_ (.A1(net212),
    .A2(_03113_),
    .B1(_02937_),
    .X(_03290_));
 nor2_1 _17690_ (.A(_02875_),
    .B(_02981_),
    .Y(_03291_));
 o21a_1 _17691_ (.A1(_03042_),
    .A2(_03291_),
    .B1(net261),
    .X(_03292_));
 or3b_1 _17692_ (.A(net218),
    .B(_02909_),
    .C_N(_03069_),
    .X(_03293_));
 a21oi_1 _17693_ (.A1(_03134_),
    .A2(_03293_),
    .B1(net267),
    .Y(_03294_));
 a311o_1 _17694_ (.A1(net267),
    .A2(_02896_),
    .A3(_02976_),
    .B1(_03294_),
    .C1(_02833_),
    .X(_03295_));
 o311a_1 _17695_ (.A1(net274),
    .A2(_03290_),
    .A3(_03292_),
    .B1(_03295_),
    .C1(net204),
    .X(_03296_));
 or3_1 _17696_ (.A(_02879_),
    .B(_02909_),
    .C(_02966_),
    .X(_03297_));
 a32o_1 _17697_ (.A1(net271),
    .A2(_03109_),
    .A3(_03136_),
    .B1(_03297_),
    .B2(_02934_),
    .X(_03298_));
 o211a_1 _17698_ (.A1(net212),
    .A2(_03069_),
    .B1(_03065_),
    .C1(net267),
    .X(_03299_));
 a31o_1 _17699_ (.A1(net261),
    .A2(_02930_),
    .A3(_02984_),
    .B1(net277),
    .X(_03300_));
 o221a_1 _17700_ (.A1(net274),
    .A2(_03298_),
    .B1(_03299_),
    .B2(_03300_),
    .C1(_02921_),
    .X(_03301_));
 o311a_4 _17701_ (.A1(net256),
    .A2(_03296_),
    .A3(_03301_),
    .B1(_03289_),
    .C1(_11361_),
    .X(_03302_));
 and2_2 _17702_ (.A(net473),
    .B(_03302_),
    .X(_03303_));
 a21o_1 _17703_ (.A1(\digitop_pav2.sec_inst.shift_in.s1.q[5] ),
    .A2(_03006_),
    .B1(_11416_),
    .X(_03304_));
 a21o_1 _17704_ (.A1(\digitop_pav2.sec_inst.shift_in.s3.q[5] ),
    .A2(net592),
    .B1(_11397_),
    .X(_03305_));
 a21o_1 _17705_ (.A1(\digitop_pav2.sec_inst.shift_in.s5.q[5] ),
    .A2(_03013_),
    .B1(net595),
    .X(_03306_));
 and4_1 _17706_ (.A(net682),
    .B(_03304_),
    .C(_03305_),
    .D(_03306_),
    .X(_03307_));
 a211o_1 _17707_ (.A1(\digitop_pav2.sec_inst.shift_in.s7.q[5] ),
    .A2(_03093_),
    .B1(_03307_),
    .C1(_11406_),
    .X(_03308_));
 and3_1 _17708_ (.A(\digitop_pav2.sec_inst.shift_in.s11.q[5] ),
    .B(net597),
    .C(_03021_),
    .X(_03309_));
 a211o_1 _17709_ (.A1(\digitop_pav2.sec_inst.shift_in.s9.q[5] ),
    .A2(_03095_),
    .B1(_03309_),
    .C1(net575),
    .X(_03310_));
 or2_1 _17710_ (.A(net1093),
    .B(net718),
    .X(_03311_));
 a31o_1 _17711_ (.A1(_03308_),
    .A2(_03310_),
    .A3(_03311_),
    .B1(net602),
    .X(_03312_));
 o211a_1 _17712_ (.A1(_08883_),
    .A2(net601),
    .B1(net535),
    .C1(_03312_),
    .X(_03313_));
 o31a_1 _17713_ (.A1(_07050_),
    .A2(net1093),
    .A3(net1017),
    .B1(net1259),
    .X(_03314_));
 o21a_2 _17714_ (.A1(_03313_),
    .A2(_03314_),
    .B1(net398),
    .X(_03315_));
 o22a_1 _17715_ (.A1(_02491_),
    .A2(_02571_),
    .B1(_02572_),
    .B2(_02490_),
    .X(_03316_));
 a22o_1 _17716_ (.A1(_02435_),
    .A2(_02485_),
    .B1(_02487_),
    .B2(_02431_),
    .X(_03317_));
 xor2_1 _17717_ (.A(_02498_),
    .B(_03317_),
    .X(_03318_));
 nand2_1 _17718_ (.A(_03316_),
    .B(_03318_),
    .Y(_03319_));
 or2_1 _17719_ (.A(_03316_),
    .B(_03318_),
    .X(_03320_));
 o21ai_1 _17720_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[13] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[13] ),
    .B1(net439),
    .Y(_03321_));
 a21oi_1 _17721_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[13] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[13] ),
    .B1(_03321_),
    .Y(_03322_));
 or2_1 _17722_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[13] ),
    .X(_03323_));
 nand2_1 _17723_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[13] ),
    .Y(_03324_));
 a31o_1 _17724_ (.A1(net427),
    .A2(_03323_),
    .A3(_03324_),
    .B1(_03322_),
    .X(_03325_));
 a311o_1 _17725_ (.A1(net470),
    .A2(_03319_),
    .A3(_03320_),
    .B1(_03325_),
    .C1(_02826_),
    .X(_03326_));
 o32a_1 _17726_ (.A1(_03303_),
    .A2(_03315_),
    .A3(_03326_),
    .B1(_02825_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[13] ),
    .X(_00409_));
 a21oi_1 _17727_ (.A1(_02910_),
    .A2(_03069_),
    .B1(net212),
    .Y(_03327_));
 a211o_1 _17728_ (.A1(net211),
    .A2(net197),
    .B1(_03327_),
    .C1(net266),
    .X(_03328_));
 o22a_1 _17729_ (.A1(_02881_),
    .A2(_02929_),
    .B1(_02991_),
    .B2(net217),
    .X(_03329_));
 o21ai_1 _17730_ (.A1(net260),
    .A2(_03329_),
    .B1(_03328_),
    .Y(_03330_));
 o32a_1 _17731_ (.A1(net219),
    .A2(_02859_),
    .A3(_02936_),
    .B1(_02908_),
    .B2(_02882_),
    .X(_03331_));
 o221a_1 _17732_ (.A1(_03071_),
    .A2(_03246_),
    .B1(_03331_),
    .B2(net262),
    .C1(net278),
    .X(_03332_));
 a211oi_1 _17733_ (.A1(net275),
    .A2(_03330_),
    .B1(_03332_),
    .C1(net203),
    .Y(_03333_));
 o211a_1 _17734_ (.A1(_02882_),
    .A2(_02908_),
    .B1(_03195_),
    .C1(net262),
    .X(_03334_));
 o31a_1 _17735_ (.A1(net217),
    .A2(_02909_),
    .A3(_02983_),
    .B1(_03072_),
    .X(_03335_));
 a21oi_1 _17736_ (.A1(_02974_),
    .A2(_03127_),
    .B1(net269),
    .Y(_03336_));
 o21ai_1 _17737_ (.A1(_03334_),
    .A2(_03335_),
    .B1(net278),
    .Y(_03337_));
 a311o_1 _17738_ (.A1(net269),
    .A2(_02928_),
    .A3(_03033_),
    .B1(_03336_),
    .C1(net279),
    .X(_03338_));
 a31o_1 _17739_ (.A1(net203),
    .A2(_03337_),
    .A3(_03338_),
    .B1(_03333_),
    .X(_03339_));
 o211a_1 _17740_ (.A1(_02877_),
    .A2(_02967_),
    .B1(_03044_),
    .C1(net259),
    .X(_03340_));
 a31o_1 _17741_ (.A1(net265),
    .A2(_02928_),
    .A3(_03032_),
    .B1(_03340_),
    .X(_03341_));
 o211a_1 _17742_ (.A1(net212),
    .A2(_02961_),
    .B1(_03195_),
    .C1(net266),
    .X(_03342_));
 a31o_1 _17743_ (.A1(net260),
    .A2(_02982_),
    .A3(_03061_),
    .B1(net273),
    .X(_03343_));
 a2bb2o_1 _17744_ (.A1_N(_03342_),
    .A2_N(_03343_),
    .B1(net273),
    .B2(_03341_),
    .X(_03344_));
 or2_1 _17745_ (.A(net194),
    .B(_02949_),
    .X(_03345_));
 o221a_1 _17746_ (.A1(net211),
    .A2(_02894_),
    .B1(net194),
    .B2(_02881_),
    .C1(net259),
    .X(_03346_));
 a31o_1 _17747_ (.A1(net270),
    .A2(_03134_),
    .A3(_03345_),
    .B1(_03346_),
    .X(_03347_));
 nor2_1 _17748_ (.A(_02899_),
    .B(_02905_),
    .Y(_03348_));
 o311a_1 _17749_ (.A1(net270),
    .A2(_03225_),
    .A3(_03348_),
    .B1(_03144_),
    .C1(net278),
    .X(_03349_));
 a211o_1 _17750_ (.A1(net275),
    .A2(_03347_),
    .B1(_03349_),
    .C1(net203),
    .X(_03350_));
 o211a_1 _17751_ (.A1(_02921_),
    .A2(_03344_),
    .B1(_03350_),
    .C1(net258),
    .X(_03351_));
 a211oi_4 _17752_ (.A1(net257),
    .A2(_03339_),
    .B1(_03351_),
    .C1(_11362_),
    .Y(_03352_));
 and2_1 _17753_ (.A(net471),
    .B(_03352_),
    .X(_03353_));
 a22o_1 _17754_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[78] ),
    .A2(net683),
    .B1(net597),
    .B2(\digitop_pav2.sec_inst.ld_r.reg96_i[62] ),
    .X(_03354_));
 a211o_1 _17755_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[94] ),
    .A2(_11417_),
    .B1(_11432_),
    .C1(_03354_),
    .X(_03355_));
 o211a_1 _17756_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[46] ),
    .A2(_11433_),
    .B1(_03355_),
    .C1(net575),
    .X(_03356_));
 or2_1 _17757_ (.A(\digitop_pav2.sec_inst.ld_r.reg96_i[14] ),
    .B(net596),
    .X(_03357_));
 o211a_1 _17758_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[30] ),
    .A2(net597),
    .B1(_11429_),
    .C1(_03357_),
    .X(_03358_));
 or4b_1 _17759_ (.A(net603),
    .B(_03356_),
    .C(_03358_),
    .D_N(net716),
    .X(_03359_));
 o221a_1 _17760_ (.A1(_08881_),
    .A2(net600),
    .B1(_10419_),
    .B2(net1089),
    .C1(net535),
    .X(_03360_));
 or3_1 _17761_ (.A(_07050_),
    .B(net1089),
    .C(net1017),
    .X(_03361_));
 a22o_1 _17762_ (.A1(_03359_),
    .A2(_03360_),
    .B1(_03361_),
    .B2(net1255),
    .X(_03362_));
 and2_2 _17763_ (.A(net398),
    .B(_03362_),
    .X(_03363_));
 or2_1 _17764_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[14] ),
    .X(_03364_));
 nand2_1 _17765_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[14] ),
    .Y(_03365_));
 or2_1 _17766_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[14] ),
    .X(_03366_));
 nand2_1 _17767_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[14] ),
    .Y(_03367_));
 a31o_1 _17768_ (.A1(net414),
    .A2(_03366_),
    .A3(_03367_),
    .B1(_02826_),
    .X(_03368_));
 a311o_1 _17769_ (.A1(net429),
    .A2(_03364_),
    .A3(_03365_),
    .B1(_03368_),
    .C1(_03363_),
    .X(_03369_));
 a22o_1 _17770_ (.A1(_02500_),
    .A2(_02585_),
    .B1(_02587_),
    .B2(_02494_),
    .X(_03370_));
 xor2_1 _17771_ (.A(_02576_),
    .B(_03370_),
    .X(_03371_));
 xnor2_1 _17772_ (.A(_02572_),
    .B(_02643_),
    .Y(_03372_));
 o21ai_1 _17773_ (.A1(_03371_),
    .A2(_03372_),
    .B1(net467),
    .Y(_03373_));
 a21oi_2 _17774_ (.A1(_03371_),
    .A2(_03372_),
    .B1(_03373_),
    .Y(_03374_));
 o32a_1 _17775_ (.A1(_03353_),
    .A2(_03369_),
    .A3(_03374_),
    .B1(_02825_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[14] ),
    .X(_00410_));
 o31a_1 _17776_ (.A1(net215),
    .A2(net210),
    .A3(net206),
    .B1(_03033_),
    .X(_03375_));
 a2111o_1 _17777_ (.A1(net220),
    .A2(_02893_),
    .B1(_02909_),
    .C1(_02870_),
    .D1(net262),
    .X(_03376_));
 o21ai_1 _17778_ (.A1(_02923_),
    .A2(_02965_),
    .B1(_03072_),
    .Y(_03377_));
 o21ai_1 _17779_ (.A1(net194),
    .A2(_02923_),
    .B1(_02905_),
    .Y(_03378_));
 o221a_1 _17780_ (.A1(_02874_),
    .A2(_02965_),
    .B1(_02989_),
    .B2(_02927_),
    .C1(net265),
    .X(_03379_));
 a21o_1 _17781_ (.A1(_02860_),
    .A2(_02981_),
    .B1(_03034_),
    .X(_03380_));
 a311o_1 _17782_ (.A1(net220),
    .A2(_02850_),
    .A3(_02873_),
    .B1(net270),
    .C1(_02902_),
    .X(_03381_));
 o32a_1 _17783_ (.A1(net217),
    .A2(_02872_),
    .A3(_02880_),
    .B1(_02980_),
    .B2(_03032_),
    .X(_03382_));
 nand2_1 _17784_ (.A(net269),
    .B(_03382_),
    .Y(_03383_));
 a31o_1 _17785_ (.A1(net219),
    .A2(net209),
    .A3(_02924_),
    .B1(_03246_),
    .X(_03384_));
 a31o_1 _17786_ (.A1(_02896_),
    .A2(_02963_),
    .A3(_02972_),
    .B1(net263),
    .X(_03385_));
 a21oi_1 _17787_ (.A1(_03384_),
    .A2(_03385_),
    .B1(net279),
    .Y(_03386_));
 a311o_1 _17788_ (.A1(net220),
    .A2(_02860_),
    .A3(_02873_),
    .B1(net269),
    .C1(_03123_),
    .X(_03387_));
 o21a_1 _17789_ (.A1(_02905_),
    .A2(_02949_),
    .B1(_02899_),
    .X(_03388_));
 o21ai_1 _17790_ (.A1(_03348_),
    .A2(_03388_),
    .B1(net269),
    .Y(_03389_));
 a311o_1 _17791_ (.A1(net279),
    .A2(_03387_),
    .A3(_03389_),
    .B1(net203),
    .C1(_03386_),
    .X(_03390_));
 o211a_1 _17792_ (.A1(net269),
    .A2(_03375_),
    .B1(_03376_),
    .C1(net278),
    .X(_03391_));
 a31o_1 _17793_ (.A1(net275),
    .A2(_03381_),
    .A3(_03383_),
    .B1(_03391_),
    .X(_03392_));
 a21oi_1 _17794_ (.A1(net203),
    .A2(_03392_),
    .B1(net258),
    .Y(_03393_));
 o311a_1 _17795_ (.A1(net270),
    .A2(_03057_),
    .A3(_03180_),
    .B1(_03377_),
    .C1(net278),
    .X(_03394_));
 o311a_1 _17796_ (.A1(net262),
    .A2(_03042_),
    .A3(_03225_),
    .B1(_03380_),
    .C1(net275),
    .X(_03395_));
 o21ai_1 _17797_ (.A1(_03394_),
    .A2(_03395_),
    .B1(net203),
    .Y(_03396_));
 a21o_1 _17798_ (.A1(net261),
    .A2(_03378_),
    .B1(_03379_),
    .X(_03397_));
 o21ba_1 _17799_ (.A1(net217),
    .A2(_03041_),
    .B1_N(_03183_),
    .X(_03398_));
 a211o_1 _17800_ (.A1(net211),
    .A2(net205),
    .B1(net265),
    .C1(_03039_),
    .X(_03399_));
 o211a_1 _17801_ (.A1(net259),
    .A2(_03398_),
    .B1(_03399_),
    .C1(net277),
    .X(_03400_));
 a211o_1 _17802_ (.A1(net273),
    .A2(_03397_),
    .B1(_03400_),
    .C1(net204),
    .X(_03401_));
 a32o_2 _17803_ (.A1(net258),
    .A2(_03396_),
    .A3(_03401_),
    .B1(_03390_),
    .B2(_03393_),
    .X(_03402_));
 and2_1 _17804_ (.A(net471),
    .B(_03402_),
    .X(_03403_));
 a22o_1 _17805_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[79] ),
    .A2(net683),
    .B1(net597),
    .B2(\digitop_pav2.sec_inst.ld_r.reg96_i[63] ),
    .X(_03404_));
 a211o_1 _17806_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[95] ),
    .A2(_11417_),
    .B1(_11432_),
    .C1(_03404_),
    .X(_03405_));
 o211a_1 _17807_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[47] ),
    .A2(_11433_),
    .B1(_03405_),
    .C1(net575),
    .X(_03406_));
 or2_1 _17808_ (.A(\digitop_pav2.sec_inst.ld_r.reg96_i[15] ),
    .B(net596),
    .X(_03407_));
 o211a_1 _17809_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[31] ),
    .A2(net597),
    .B1(_11429_),
    .C1(_03407_),
    .X(_03408_));
 or4b_1 _17810_ (.A(net603),
    .B(_03406_),
    .C(_03408_),
    .D_N(net717),
    .X(_03409_));
 o221a_1 _17811_ (.A1(_08880_),
    .A2(net600),
    .B1(_10419_),
    .B2(net1086),
    .C1(net534),
    .X(_03410_));
 a22o_1 _17812_ (.A1(net1086),
    .A2(_02414_),
    .B1(_03409_),
    .B2(_03410_),
    .X(_03411_));
 and2_2 _17813_ (.A(net398),
    .B(_03411_),
    .X(_03412_));
 o21ai_1 _17814_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[15] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[15] ),
    .B1(net429),
    .Y(_03413_));
 a21oi_1 _17815_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[15] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[15] ),
    .B1(_03413_),
    .Y(_03414_));
 xor2_1 _17816_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[15] ),
    .X(_03415_));
 a2111o_1 _17817_ (.A1(net415),
    .A2(_03415_),
    .B1(_03414_),
    .C1(_03412_),
    .D1(_02826_),
    .X(_03416_));
 a22o_1 _17818_ (.A1(_02580_),
    .A2(_02634_),
    .B1(_02636_),
    .B2(_02579_),
    .X(_03417_));
 xnor2_1 _17819_ (.A(_11456_),
    .B(_03417_),
    .Y(_03418_));
 xnor2_1 _17820_ (.A(_11463_),
    .B(_02643_),
    .Y(_03419_));
 o21ai_1 _17821_ (.A1(_03418_),
    .A2(_03419_),
    .B1(net467),
    .Y(_03420_));
 a21oi_2 _17822_ (.A1(_03418_),
    .A2(_03419_),
    .B1(_03420_),
    .Y(_03421_));
 o32a_1 _17823_ (.A1(_03403_),
    .A2(_03416_),
    .A3(_03421_),
    .B1(_02825_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[15] ),
    .X(_00411_));
 nand2_4 _17824_ (.A(net468),
    .B(_11446_),
    .Y(_03422_));
 o21ai_2 _17825_ (.A1(_11191_),
    .A2(_11193_),
    .B1(_03422_),
    .Y(_03423_));
 and2_1 _17826_ (.A(net417),
    .B(net173),
    .X(_03424_));
 nand2_2 _17827_ (.A(net417),
    .B(net173),
    .Y(_03425_));
 a22o_1 _17828_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[4] ),
    .A2(net358),
    .B1(_11214_),
    .B2(_07517_),
    .X(_03426_));
 nand2_2 _17829_ (.A(_10743_),
    .B(_03426_),
    .Y(_03427_));
 and3b_2 _17830_ (.A_N(_03423_),
    .B(_03425_),
    .C(_03427_),
    .X(_03428_));
 or3b_4 _17831_ (.A(_03423_),
    .B(_03424_),
    .C_N(_03427_),
    .X(_03429_));
 nand2_1 _17832_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[8] ),
    .Y(_03430_));
 or2_1 _17833_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[8] ),
    .X(_03431_));
 a311o_1 _17834_ (.A1(net402),
    .A2(_03430_),
    .A3(_03431_),
    .B1(_03026_),
    .C1(_03429_),
    .X(_03432_));
 a22o_1 _17835_ (.A1(_11471_),
    .A2(_02206_),
    .B1(_02207_),
    .B2(_11470_),
    .X(_03433_));
 xnor2_2 _17836_ (.A(_11456_),
    .B(_03433_),
    .Y(_03434_));
 o21ai_1 _17837_ (.A1(_02754_),
    .A2(_03434_),
    .B1(net466),
    .Y(_03435_));
 a21oi_4 _17838_ (.A1(_02754_),
    .A2(_03434_),
    .B1(_03435_),
    .Y(_03436_));
 o32a_1 _17839_ (.A1(_02996_),
    .A2(_03432_),
    .A3(_03436_),
    .B1(_03428_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[8] ),
    .X(_00412_));
 nand2_1 _17840_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[9] ),
    .Y(_03437_));
 or2_1 _17841_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[9] ),
    .X(_03438_));
 a311o_1 _17842_ (.A1(net399),
    .A2(_03437_),
    .A3(_03438_),
    .B1(_03101_),
    .C1(_03429_),
    .X(_03439_));
 xnor2_1 _17843_ (.A(_02196_),
    .B(_02290_),
    .Y(_03440_));
 xnor2_1 _17844_ (.A(_11458_),
    .B(_03440_),
    .Y(_03441_));
 xnor2_1 _17845_ (.A(_02201_),
    .B(_02754_),
    .Y(_03442_));
 o21ai_1 _17846_ (.A1(_03441_),
    .A2(_03442_),
    .B1(net466),
    .Y(_03443_));
 a21oi_2 _17847_ (.A1(_03441_),
    .A2(_03442_),
    .B1(_03443_),
    .Y(_03444_));
 o32a_1 _17848_ (.A1(_03082_),
    .A2(_03439_),
    .A3(_03444_),
    .B1(_03428_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[9] ),
    .X(_00413_));
 xor2_1 _17849_ (.A(_02212_),
    .B(_02299_),
    .X(_03445_));
 a22o_1 _17850_ (.A1(_02202_),
    .A2(_02294_),
    .B1(_02295_),
    .B2(_02200_),
    .X(_03446_));
 xnor2_1 _17851_ (.A(_03445_),
    .B(_03446_),
    .Y(_03447_));
 a21boi_1 _17852_ (.A1(_02357_),
    .A2(_03447_),
    .B1_N(net466),
    .Y(_03448_));
 o21a_1 _17853_ (.A1(_02357_),
    .A2(_03447_),
    .B1(_03448_),
    .X(_03449_));
 or2_1 _17854_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[10] ),
    .X(_03450_));
 nand2_1 _17855_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[10] ),
    .Y(_03451_));
 a311o_1 _17856_ (.A1(net400),
    .A2(_03450_),
    .A3(_03451_),
    .B1(_03162_),
    .C1(_03429_),
    .X(_03452_));
 o32a_1 _17857_ (.A1(_03150_),
    .A2(_03449_),
    .A3(_03452_),
    .B1(_03428_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[10] ),
    .X(_00414_));
 nand2_1 _17858_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[11] ),
    .Y(_03453_));
 or2_1 _17859_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[11] ),
    .X(_03454_));
 a311o_1 _17860_ (.A1(net402),
    .A2(_03453_),
    .A3(_03454_),
    .B1(_03217_),
    .C1(_03429_),
    .X(_03455_));
 o22a_1 _17861_ (.A1(_02368_),
    .A2(_02427_),
    .B1(_02428_),
    .B2(_02367_),
    .X(_03456_));
 xor2_1 _17862_ (.A(_11456_),
    .B(_02284_),
    .X(_03457_));
 xnor2_1 _17863_ (.A(_03456_),
    .B(_03457_),
    .Y(_03458_));
 xnor2_1 _17864_ (.A(_02362_),
    .B(_02774_),
    .Y(_03459_));
 o21ai_1 _17865_ (.A1(_03458_),
    .A2(_03459_),
    .B1(net468),
    .Y(_03460_));
 a21oi_2 _17866_ (.A1(_03458_),
    .A2(_03459_),
    .B1(_03460_),
    .Y(_03461_));
 o32a_1 _17867_ (.A1(_03202_),
    .A2(_03455_),
    .A3(_03461_),
    .B1(_03428_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[11] ),
    .X(_00415_));
 nand2_1 _17868_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[12] ),
    .Y(_03462_));
 or2_1 _17869_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[12] ),
    .X(_03463_));
 a311o_1 _17870_ (.A1(net402),
    .A2(_03462_),
    .A3(_03463_),
    .B1(_03269_),
    .C1(_03429_),
    .X(_03464_));
 xor2_1 _17871_ (.A(_02435_),
    .B(_02491_),
    .X(_03465_));
 xnor2_1 _17872_ (.A(_02375_),
    .B(_03465_),
    .Y(_03466_));
 xnor2_1 _17873_ (.A(_02434_),
    .B(_02783_),
    .Y(_03467_));
 o21ai_1 _17874_ (.A1(_03466_),
    .A2(_03467_),
    .B1(net469),
    .Y(_03468_));
 a21oi_2 _17875_ (.A1(_03466_),
    .A2(_03467_),
    .B1(_03468_),
    .Y(_03469_));
 o32a_1 _17876_ (.A1(_03255_),
    .A2(_03464_),
    .A3(_03469_),
    .B1(_03428_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[12] ),
    .X(_00416_));
 nand2_1 _17877_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[13] ),
    .Y(_03470_));
 or2_1 _17878_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[13] ),
    .X(_03471_));
 a311o_1 _17879_ (.A1(net402),
    .A2(_03470_),
    .A3(_03471_),
    .B1(_03315_),
    .C1(_03429_),
    .X(_03472_));
 mux2_1 _17880_ (.A0(_02497_),
    .A1(_02498_),
    .S(_02434_),
    .X(_03473_));
 xnor2_1 _17881_ (.A(_02439_),
    .B(_02572_),
    .Y(_03474_));
 xnor2_1 _17882_ (.A(_02499_),
    .B(_03474_),
    .Y(_03475_));
 o21ai_1 _17883_ (.A1(_03473_),
    .A2(_03475_),
    .B1(net469),
    .Y(_03476_));
 a21oi_2 _17884_ (.A1(_03473_),
    .A2(_03475_),
    .B1(_03476_),
    .Y(_03477_));
 o32a_1 _17885_ (.A1(_03303_),
    .A2(_03472_),
    .A3(_03477_),
    .B1(_03428_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[13] ),
    .X(_00417_));
 xnor2_1 _17886_ (.A(_02498_),
    .B(_02576_),
    .Y(_03478_));
 xnor2_1 _17887_ (.A(_02486_),
    .B(_02580_),
    .Y(_03479_));
 xnor2_1 _17888_ (.A(_02643_),
    .B(_03479_),
    .Y(_03480_));
 xnor2_1 _17889_ (.A(_03478_),
    .B(_03480_),
    .Y(_03481_));
 a21o_1 _17890_ (.A1(net466),
    .A2(_03481_),
    .B1(_03353_),
    .X(_03482_));
 or2_1 _17891_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[14] ),
    .X(_03483_));
 nand2_1 _17892_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[14] ),
    .Y(_03484_));
 a31o_1 _17893_ (.A1(net399),
    .A2(_03483_),
    .A3(_03484_),
    .B1(_03429_),
    .X(_03485_));
 o32a_1 _17894_ (.A1(_03363_),
    .A2(_03482_),
    .A3(_03485_),
    .B1(_03428_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[14] ),
    .X(_00418_));
 a22o_1 _17895_ (.A1(_11462_),
    .A2(_02585_),
    .B1(_02587_),
    .B2(_11461_),
    .X(_03486_));
 xnor2_1 _17896_ (.A(_02644_),
    .B(_03486_),
    .Y(_03487_));
 mux2_1 _17897_ (.A0(_02575_),
    .A1(_02576_),
    .S(_02635_),
    .X(_03488_));
 o21ai_1 _17898_ (.A1(_03487_),
    .A2(_03488_),
    .B1(net467),
    .Y(_03489_));
 a21oi_1 _17899_ (.A1(_03487_),
    .A2(_03488_),
    .B1(_03489_),
    .Y(_03490_));
 or2_1 _17900_ (.A(_03403_),
    .B(_03490_),
    .X(_03491_));
 or2_1 _17901_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[15] ),
    .X(_03492_));
 nand2_1 _17902_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[15] ),
    .Y(_03493_));
 a31o_1 _17903_ (.A1(net399),
    .A2(_03492_),
    .A3(_03493_),
    .B1(_03429_),
    .X(_03494_));
 o32a_1 _17904_ (.A1(_03412_),
    .A2(_03491_),
    .A3(_03494_),
    .B1(_03428_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[15] ),
    .X(_00419_));
 o22a_2 _17905_ (.A1(_11192_),
    .A2(net357),
    .B1(net389),
    .B2(_07516_),
    .X(_03495_));
 and3_2 _17906_ (.A(_11198_),
    .B(_02824_),
    .C(_03495_),
    .X(_03496_));
 nand3_4 _17907_ (.A(_11198_),
    .B(_02824_),
    .C(_03495_),
    .Y(_03497_));
 o21ai_1 _17908_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[8] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[8] ),
    .B1(net438),
    .Y(_03498_));
 a21oi_1 _17909_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[8] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[8] ),
    .B1(_03498_),
    .Y(_03499_));
 xor2_1 _17910_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[8] ),
    .X(_03500_));
 a211o_1 _17911_ (.A1(net425),
    .A2(_03500_),
    .B1(_03499_),
    .C1(_03497_),
    .X(_03501_));
 o32a_1 _17912_ (.A1(_02996_),
    .A2(_03031_),
    .A3(_03501_),
    .B1(_03496_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[8] ),
    .X(_00420_));
 o21ai_1 _17913_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[9] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[9] ),
    .B1(net429),
    .Y(_03502_));
 a21oi_1 _17914_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[9] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[9] ),
    .B1(_03502_),
    .Y(_03503_));
 or2_1 _17915_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[9] ),
    .X(_03504_));
 nand2_1 _17916_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[9] ),
    .Y(_03505_));
 a31o_1 _17917_ (.A1(net414),
    .A2(_03504_),
    .A3(_03505_),
    .B1(_03503_),
    .X(_03506_));
 or4b_1 _17918_ (.A(_03082_),
    .B(_03497_),
    .C(_03506_),
    .D_N(_03106_),
    .X(_03507_));
 o22a_1 _17919_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[9] ),
    .A2(_03496_),
    .B1(_03507_),
    .B2(_03101_),
    .X(_00421_));
 or2_1 _17920_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[10] ),
    .X(_03508_));
 nand2_1 _17921_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[10] ),
    .Y(_03509_));
 or2_1 _17922_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[10] ),
    .X(_03510_));
 nand2_1 _17923_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[10] ),
    .Y(_03511_));
 a311o_1 _17924_ (.A1(net416),
    .A2(_03508_),
    .A3(_03509_),
    .B1(_03162_),
    .C1(_03497_),
    .X(_03512_));
 a31o_1 _17925_ (.A1(net431),
    .A2(_03510_),
    .A3(_03511_),
    .B1(_03512_),
    .X(_03513_));
 o32a_1 _17926_ (.A1(_03150_),
    .A2(_03171_),
    .A3(_03513_),
    .B1(_03496_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ),
    .X(_00422_));
 o21ai_1 _17927_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[11] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[11] ),
    .B1(net438),
    .Y(_03514_));
 a21oi_1 _17928_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[11] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[11] ),
    .B1(_03514_),
    .Y(_03515_));
 xor2_1 _17929_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[11] ),
    .X(_03516_));
 a2111o_1 _17930_ (.A1(net425),
    .A2(_03516_),
    .B1(_03515_),
    .C1(_03497_),
    .D1(_03217_),
    .X(_03517_));
 o32a_1 _17931_ (.A1(_03202_),
    .A2(_03223_),
    .A3(_03517_),
    .B1(_03496_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[11] ),
    .X(_00423_));
 o21ai_1 _17932_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[12] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[12] ),
    .B1(net438),
    .Y(_03518_));
 a21oi_1 _17933_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[12] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[12] ),
    .B1(_03518_),
    .Y(_03519_));
 xor2_1 _17934_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[12] ),
    .X(_03520_));
 a2111o_1 _17935_ (.A1(net425),
    .A2(_03520_),
    .B1(_03519_),
    .C1(_03497_),
    .D1(_03269_),
    .X(_03521_));
 o32a_1 _17936_ (.A1(_03255_),
    .A2(_03274_),
    .A3(_03521_),
    .B1(_03496_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[12] ),
    .X(_00424_));
 o21ai_1 _17937_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[13] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[13] ),
    .B1(net438),
    .Y(_03522_));
 a21oi_1 _17938_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[13] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[13] ),
    .B1(_03522_),
    .Y(_03523_));
 xor2_1 _17939_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[13] ),
    .X(_03524_));
 a211o_1 _17940_ (.A1(net425),
    .A2(_03524_),
    .B1(_03523_),
    .C1(_03497_),
    .X(_03525_));
 a31o_1 _17941_ (.A1(net470),
    .A2(_03319_),
    .A3(_03320_),
    .B1(_03315_),
    .X(_03526_));
 o32a_1 _17942_ (.A1(_03303_),
    .A2(_03525_),
    .A3(_03526_),
    .B1(_03496_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[13] ),
    .X(_00425_));
 xor2_1 _17943_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[14] ),
    .X(_03527_));
 o21ai_1 _17944_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[14] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[14] ),
    .B1(net429),
    .Y(_03528_));
 a21oi_1 _17945_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[14] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[14] ),
    .B1(_03528_),
    .Y(_03529_));
 a2111o_1 _17946_ (.A1(net414),
    .A2(_03527_),
    .B1(_03529_),
    .C1(_03363_),
    .D1(_03497_),
    .X(_03530_));
 o32a_1 _17947_ (.A1(_03353_),
    .A2(_03374_),
    .A3(_03530_),
    .B1(_03496_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[14] ),
    .X(_00426_));
 o21ai_1 _17948_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[15] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[15] ),
    .B1(net430),
    .Y(_03531_));
 a21oi_1 _17949_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[15] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[15] ),
    .B1(_03531_),
    .Y(_03532_));
 xor2_1 _17950_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[15] ),
    .X(_03533_));
 a2111o_1 _17951_ (.A1(net414),
    .A2(_03533_),
    .B1(_03532_),
    .C1(_03497_),
    .D1(_03412_),
    .X(_03534_));
 o32a_1 _17952_ (.A1(_03403_),
    .A2(_03421_),
    .A3(_03534_),
    .B1(_03496_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[15] ),
    .X(_00427_));
 o2bb2a_1 _17953_ (.A1_N(_07517_),
    .A2_N(_11202_),
    .B1(net389),
    .B2(_11192_),
    .X(_03535_));
 a22o_1 _17954_ (.A1(_07517_),
    .A2(_11202_),
    .B1(_11216_),
    .B2(_11191_),
    .X(_03536_));
 and3b_4 _17955_ (.A_N(_03423_),
    .B(_03535_),
    .C(_02735_),
    .X(_03537_));
 or3b_4 _17956_ (.A(_03423_),
    .B(_03536_),
    .C_N(_02735_),
    .X(_03538_));
 xor2_1 _17957_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[0] ),
    .X(_03539_));
 o21ai_1 _17958_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[0] ),
    .B1(net433),
    .Y(_03540_));
 a21oi_1 _17959_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[0] ),
    .B1(_03540_),
    .Y(_03541_));
 a211o_1 _17960_ (.A1(net420),
    .A2(_03539_),
    .B1(_03541_),
    .C1(_03538_),
    .X(_03542_));
 o32a_1 _17961_ (.A1(_11393_),
    .A2(_02747_),
    .A3(_03542_),
    .B1(_03537_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[0] ),
    .X(_00428_));
 o21ai_1 _17962_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[1] ),
    .B1(net434),
    .Y(_03543_));
 a21oi_1 _17963_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[1] ),
    .B1(_03543_),
    .Y(_03544_));
 xor2_1 _17964_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[1] ),
    .X(_03545_));
 a211o_1 _17965_ (.A1(net418),
    .A2(_03545_),
    .B1(_03544_),
    .C1(_03538_),
    .X(_03546_));
 o32a_1 _17966_ (.A1(_02182_),
    .A2(_02758_),
    .A3(_03546_),
    .B1(_03537_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[1] ),
    .X(_00429_));
 o21ai_1 _17967_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[2] ),
    .B1(net435),
    .Y(_03547_));
 a21oi_1 _17968_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[2] ),
    .B1(_03547_),
    .Y(_03548_));
 xor2_1 _17969_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[2] ),
    .X(_03549_));
 a2111o_1 _17970_ (.A1(net421),
    .A2(_03549_),
    .B1(_03548_),
    .C1(_03538_),
    .D1(_02280_),
    .X(_03550_));
 o32a_1 _17971_ (.A1(_02265_),
    .A2(_02767_),
    .A3(_03550_),
    .B1(_03537_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[2] ),
    .X(_00430_));
 or2_1 _17972_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[3] ),
    .X(_03551_));
 nand2_1 _17973_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[3] ),
    .Y(_03552_));
 or2_1 _17974_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[3] ),
    .X(_03553_));
 nand2_1 _17975_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[3] ),
    .Y(_03554_));
 a311o_1 _17976_ (.A1(net436),
    .A2(_03553_),
    .A3(_03554_),
    .B1(_02354_),
    .C1(_03538_),
    .X(_03555_));
 a31o_1 _17977_ (.A1(net422),
    .A2(_03551_),
    .A3(_03552_),
    .B1(_03555_),
    .X(_03556_));
 o32a_1 _17978_ (.A1(_02339_),
    .A2(_02779_),
    .A3(_03556_),
    .B1(_03537_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[3] ),
    .X(_00431_));
 o21ai_1 _17979_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[4] ),
    .B1(net437),
    .Y(_03557_));
 a21oi_1 _17980_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[4] ),
    .B1(_03557_),
    .Y(_03558_));
 xor2_1 _17981_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[4] ),
    .X(_03559_));
 a2111o_1 _17982_ (.A1(net423),
    .A2(_03559_),
    .B1(_03558_),
    .C1(_03538_),
    .D1(_02423_),
    .X(_03560_));
 o32a_1 _17983_ (.A1(_02413_),
    .A2(_02788_),
    .A3(_03560_),
    .B1(_03537_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[4] ),
    .X(_00432_));
 o21ai_1 _17984_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[5] ),
    .B1(net437),
    .Y(_03561_));
 a21oi_1 _17985_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[5] ),
    .B1(_03561_),
    .Y(_03562_));
 or2_1 _17986_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[5] ),
    .X(_03563_));
 nand2_1 _17987_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[5] ),
    .Y(_03564_));
 a31o_1 _17988_ (.A1(net423),
    .A2(_03563_),
    .A3(_03564_),
    .B1(_03562_),
    .X(_03565_));
 or4_1 _17989_ (.A(_02511_),
    .B(_02794_),
    .C(_03538_),
    .D(_03565_),
    .X(_03566_));
 o22a_1 _17990_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[5] ),
    .A2(_03537_),
    .B1(_03566_),
    .B2(_02482_),
    .X(_00433_));
 or2_1 _17991_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[6] ),
    .X(_03567_));
 nand2_1 _17992_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[6] ),
    .Y(_03568_));
 or2_1 _17993_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[6] ),
    .X(_03569_));
 nand2_1 _17994_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[6] ),
    .Y(_03570_));
 a311o_1 _17995_ (.A1(net432),
    .A2(_03567_),
    .A3(_03568_),
    .B1(_02562_),
    .C1(_02811_),
    .X(_03571_));
 a31o_1 _17996_ (.A1(net418),
    .A2(_03569_),
    .A3(_03570_),
    .B1(_03538_),
    .X(_03572_));
 o32a_1 _17997_ (.A1(_02552_),
    .A2(_03571_),
    .A3(_03572_),
    .B1(_03537_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[6] ),
    .X(_00434_));
 o21ai_1 _17998_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[7] ),
    .B1(net415),
    .Y(_03573_));
 a21oi_1 _17999_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[7] ),
    .B1(_03573_),
    .Y(_03574_));
 or2_1 _18000_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[7] ),
    .X(_03575_));
 nand2_1 _18001_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[7] ),
    .Y(_03576_));
 a311o_1 _18002_ (.A1(net430),
    .A2(_03575_),
    .A3(_03576_),
    .B1(_03538_),
    .C1(_03574_),
    .X(_03577_));
 o32a_1 _18003_ (.A1(_02616_),
    .A2(_02821_),
    .A3(_03577_),
    .B1(_03537_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[7] ),
    .X(_00435_));
 or2_1 _18004_ (.A(_07516_),
    .B(net354),
    .X(_03578_));
 a31o_2 _18005_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[4] ),
    .A2(_10743_),
    .A3(net364),
    .B1(_11193_),
    .X(_03579_));
 and4_4 _18006_ (.A(_02735_),
    .B(_02823_),
    .C(_03578_),
    .D(_03579_),
    .X(_03580_));
 nand4_4 _18007_ (.A(_02735_),
    .B(_02823_),
    .C(_03578_),
    .D(_03579_),
    .Y(_03581_));
 xor2_1 _18008_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[0] ),
    .X(_03582_));
 o21ai_1 _18009_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[0] ),
    .B1(net433),
    .Y(_03583_));
 a21oi_1 _18010_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[0] ),
    .B1(_03583_),
    .Y(_03584_));
 a211o_1 _18011_ (.A1(net419),
    .A2(_03582_),
    .B1(_03584_),
    .C1(_03581_),
    .X(_03585_));
 o32a_1 _18012_ (.A1(_11393_),
    .A2(_02747_),
    .A3(_03585_),
    .B1(_03580_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[0] ),
    .X(_00436_));
 o21ai_1 _18013_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[1] ),
    .B1(net432),
    .Y(_03586_));
 a21oi_1 _18014_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[1] ),
    .B1(_03586_),
    .Y(_03587_));
 xor2_1 _18015_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[1] ),
    .X(_03588_));
 a211o_1 _18016_ (.A1(net418),
    .A2(_03588_),
    .B1(_03587_),
    .C1(_03581_),
    .X(_03589_));
 o32a_1 _18017_ (.A1(_02182_),
    .A2(_02758_),
    .A3(_03589_),
    .B1(_03580_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[1] ),
    .X(_00437_));
 or2_1 _18018_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[2] ),
    .X(_03590_));
 nand2_1 _18019_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[2] ),
    .Y(_03591_));
 or2_1 _18020_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[2] ),
    .X(_03592_));
 nand2_1 _18021_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[2] ),
    .Y(_03593_));
 a31o_1 _18022_ (.A1(net421),
    .A2(_03592_),
    .A3(_03593_),
    .B1(_03581_),
    .X(_03594_));
 a311o_1 _18023_ (.A1(net435),
    .A2(_03590_),
    .A3(_03591_),
    .B1(_03594_),
    .C1(_02280_),
    .X(_03595_));
 o32a_1 _18024_ (.A1(_02265_),
    .A2(_02767_),
    .A3(_03595_),
    .B1(_03580_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[2] ),
    .X(_00438_));
 o21ai_1 _18025_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[3] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[3] ),
    .B1(net419),
    .Y(_03596_));
 a21oi_1 _18026_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[3] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[3] ),
    .B1(_03596_),
    .Y(_03597_));
 xor2_1 _18027_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[3] ),
    .X(_03598_));
 a2111o_1 _18028_ (.A1(net436),
    .A2(_03598_),
    .B1(_03597_),
    .C1(_03581_),
    .D1(_02354_),
    .X(_03599_));
 o32a_1 _18029_ (.A1(_02339_),
    .A2(_02779_),
    .A3(_03599_),
    .B1(_03580_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[3] ),
    .X(_00439_));
 o21ai_1 _18030_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[4] ),
    .B1(net437),
    .Y(_03600_));
 a21oi_1 _18031_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[4] ),
    .B1(_03600_),
    .Y(_03601_));
 xor2_1 _18032_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[4] ),
    .X(_03602_));
 a2111o_1 _18033_ (.A1(net424),
    .A2(_03602_),
    .B1(_03601_),
    .C1(_03581_),
    .D1(_02423_),
    .X(_03603_));
 o32a_1 _18034_ (.A1(_02413_),
    .A2(_02788_),
    .A3(_03603_),
    .B1(_03580_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[4] ),
    .X(_00440_));
 o21ai_1 _18035_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[5] ),
    .B1(net437),
    .Y(_03604_));
 a21oi_1 _18036_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[5] ),
    .B1(_03604_),
    .Y(_03605_));
 or2_1 _18037_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[5] ),
    .X(_03606_));
 nand2_1 _18038_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[5] ),
    .Y(_03607_));
 a31o_1 _18039_ (.A1(net422),
    .A2(_03606_),
    .A3(_03607_),
    .B1(_03605_),
    .X(_03608_));
 or4_1 _18040_ (.A(_02511_),
    .B(_02794_),
    .C(_03581_),
    .D(_03608_),
    .X(_03609_));
 o22a_1 _18041_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[5] ),
    .A2(_03580_),
    .B1(_03609_),
    .B2(_02482_),
    .X(_00441_));
 o21ai_1 _18042_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[6] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[6] ),
    .B1(net432),
    .Y(_03610_));
 a21oi_1 _18043_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[6] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[6] ),
    .B1(_03610_),
    .Y(_03611_));
 xor2_1 _18044_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[6] ),
    .X(_03612_));
 a2111o_1 _18045_ (.A1(net418),
    .A2(_03612_),
    .B1(_03611_),
    .C1(_03581_),
    .D1(_02562_),
    .X(_03613_));
 o32a_1 _18046_ (.A1(_02552_),
    .A2(_02811_),
    .A3(_03613_),
    .B1(_03580_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[6] ),
    .X(_00442_));
 or2_1 _18047_ (.A(_02616_),
    .B(_02821_),
    .X(_03614_));
 xor2_1 _18048_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[7] ),
    .X(_03615_));
 o21ai_1 _18049_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[7] ),
    .B1(net435),
    .Y(_03616_));
 a21oi_1 _18050_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[7] ),
    .B1(_03616_),
    .Y(_03617_));
 a211o_1 _18051_ (.A1(net421),
    .A2(_03615_),
    .B1(_03617_),
    .C1(_03581_),
    .X(_03618_));
 o22a_1 _18052_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ),
    .A2(_03580_),
    .B1(_03614_),
    .B2(_03618_),
    .X(_00443_));
 o22a_2 _18053_ (.A1(_07516_),
    .A2(net391),
    .B1(net355),
    .B2(_11192_),
    .X(_03619_));
 and3_2 _18054_ (.A(_02824_),
    .B(_03422_),
    .C(_03619_),
    .X(_03620_));
 nand3_4 _18055_ (.A(_02824_),
    .B(_03422_),
    .C(_03619_),
    .Y(_03621_));
 o21ai_1 _18056_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[8] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[8] ),
    .B1(net431),
    .Y(_03622_));
 a21oi_1 _18057_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[8] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[8] ),
    .B1(_03622_),
    .Y(_03623_));
 xor2_1 _18058_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[8] ),
    .X(_03624_));
 a211o_1 _18059_ (.A1(net416),
    .A2(_03624_),
    .B1(_03623_),
    .C1(_03621_),
    .X(_03625_));
 o32a_1 _18060_ (.A1(_02996_),
    .A2(_03031_),
    .A3(_03625_),
    .B1(_03620_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[8] ),
    .X(_00444_));
 o21ai_1 _18061_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[9] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[9] ),
    .B1(net429),
    .Y(_03626_));
 a21oi_1 _18062_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[9] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[9] ),
    .B1(_03626_),
    .Y(_03627_));
 or2_1 _18063_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[9] ),
    .X(_03628_));
 nand2_1 _18064_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[9] ),
    .Y(_03629_));
 a31o_1 _18065_ (.A1(net414),
    .A2(_03628_),
    .A3(_03629_),
    .B1(_03627_),
    .X(_03630_));
 or4b_1 _18066_ (.A(_03082_),
    .B(_03621_),
    .C(_03630_),
    .D_N(_03106_),
    .X(_03631_));
 o22a_1 _18067_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[9] ),
    .A2(_03620_),
    .B1(_03631_),
    .B2(_03101_),
    .X(_00445_));
 or2_1 _18068_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[10] ),
    .X(_03632_));
 nand2_1 _18069_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[10] ),
    .Y(_03633_));
 or2_1 _18070_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[10] ),
    .X(_03634_));
 nand2_1 _18071_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[10] ),
    .Y(_03635_));
 a311o_1 _18072_ (.A1(net416),
    .A2(_03632_),
    .A3(_03633_),
    .B1(_03162_),
    .C1(_03621_),
    .X(_03636_));
 a31o_1 _18073_ (.A1(net431),
    .A2(_03634_),
    .A3(_03635_),
    .B1(_03636_),
    .X(_03637_));
 o32a_1 _18074_ (.A1(_03150_),
    .A2(_03171_),
    .A3(_03637_),
    .B1(_03620_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[10] ),
    .X(_00446_));
 o21ai_1 _18075_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[11] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[11] ),
    .B1(net438),
    .Y(_03638_));
 a21oi_1 _18076_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[11] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[11] ),
    .B1(_03638_),
    .Y(_03639_));
 xor2_1 _18077_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[11] ),
    .X(_03640_));
 a2111o_1 _18078_ (.A1(net425),
    .A2(_03640_),
    .B1(_03639_),
    .C1(_03621_),
    .D1(_03217_),
    .X(_03641_));
 o32a_1 _18079_ (.A1(_03202_),
    .A2(_03223_),
    .A3(_03641_),
    .B1(_03620_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[11] ),
    .X(_00447_));
 o21ai_1 _18080_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[12] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[12] ),
    .B1(net431),
    .Y(_03642_));
 a21oi_1 _18081_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[12] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[12] ),
    .B1(_03642_),
    .Y(_03643_));
 xor2_1 _18082_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[12] ),
    .X(_03644_));
 a2111o_1 _18083_ (.A1(net416),
    .A2(_03644_),
    .B1(_03643_),
    .C1(_03621_),
    .D1(_03269_),
    .X(_03645_));
 o32a_1 _18084_ (.A1(_03255_),
    .A2(_03274_),
    .A3(_03645_),
    .B1(_03620_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[12] ),
    .X(_00448_));
 o21ai_1 _18085_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[13] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[13] ),
    .B1(net438),
    .Y(_03646_));
 a21oi_1 _18086_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[13] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[13] ),
    .B1(_03646_),
    .Y(_03647_));
 xor2_1 _18087_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[13] ),
    .X(_03648_));
 a211o_1 _18088_ (.A1(net425),
    .A2(_03648_),
    .B1(_03647_),
    .C1(_03621_),
    .X(_03649_));
 o32a_1 _18089_ (.A1(_03303_),
    .A2(_03526_),
    .A3(_03649_),
    .B1(_03620_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[13] ),
    .X(_00449_));
 or2_1 _18090_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[14] ),
    .X(_03650_));
 nand2_1 _18091_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[14] ),
    .Y(_03651_));
 o21ai_1 _18092_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[14] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[14] ),
    .B1(net429),
    .Y(_03652_));
 a21oi_1 _18093_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[14] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[14] ),
    .B1(_03652_),
    .Y(_03653_));
 a31o_1 _18094_ (.A1(net414),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_03653_),
    .X(_03654_));
 or3_1 _18095_ (.A(_03363_),
    .B(_03621_),
    .C(_03654_),
    .X(_03655_));
 o32a_1 _18096_ (.A1(_03353_),
    .A2(_03374_),
    .A3(_03655_),
    .B1(_03620_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[14] ),
    .X(_00450_));
 o21ai_1 _18097_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[15] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[15] ),
    .B1(net429),
    .Y(_03656_));
 a21oi_1 _18098_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[15] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[15] ),
    .B1(_03656_),
    .Y(_03657_));
 xor2_1 _18099_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[15] ),
    .X(_03658_));
 a2111o_1 _18100_ (.A1(net414),
    .A2(_03658_),
    .B1(_03657_),
    .C1(_03621_),
    .D1(_03412_),
    .X(_03659_));
 o32a_1 _18101_ (.A1(_03403_),
    .A2(_03421_),
    .A3(_03659_),
    .B1(_03620_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[15] ),
    .X(_00451_));
 or3b_1 _18102_ (.A(_07832_),
    .B(net1326),
    .C_N(\digitop_pav2.boot_inst.boot_proc0.proc_stage[1] ),
    .X(_03660_));
 mux2_1 _18103_ (.A0(net1134),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[0] ),
    .S(net1312),
    .X(_00452_));
 mux2_1 _18104_ (.A0(net1133),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[1] ),
    .S(net1312),
    .X(_00453_));
 mux2_1 _18105_ (.A0(net1127),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[2] ),
    .S(net1312),
    .X(_00454_));
 mux2_1 _18106_ (.A0(net1124),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[3] ),
    .S(net1312),
    .X(_00455_));
 mux2_1 _18107_ (.A0(net1121),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[4] ),
    .S(net1312),
    .X(_00456_));
 mux2_1 _18108_ (.A0(net1118),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[5] ),
    .S(net1312),
    .X(_00457_));
 mux2_1 _18109_ (.A0(net1116),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[6] ),
    .S(net1313),
    .X(_00458_));
 mux2_1 _18110_ (.A0(net1113),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[7] ),
    .S(net1312),
    .X(_00459_));
 mux2_1 _18111_ (.A0(net1107),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[8] ),
    .S(net1313),
    .X(_00460_));
 mux2_1 _18112_ (.A0(net1105),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[9] ),
    .S(net1313),
    .X(_00461_));
 mux2_1 _18113_ (.A0(net1100),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[10] ),
    .S(net1313),
    .X(_00462_));
 mux2_1 _18114_ (.A0(net1096),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[11] ),
    .S(net1313),
    .X(_00463_));
 mux2_1 _18115_ (.A0(net1095),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[12] ),
    .S(net1313),
    .X(_00464_));
 mux2_1 _18116_ (.A0(net1092),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[13] ),
    .S(net1312),
    .X(_00465_));
 mux2_1 _18117_ (.A0(net1087),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[14] ),
    .S(net1312),
    .X(_00466_));
 mux2_1 _18118_ (.A0(net1085),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[15] ),
    .S(net1312),
    .X(_00467_));
 nor3_1 _18119_ (.A(net1248),
    .B(net818),
    .C(net1712),
    .Y(_03661_));
 or3_2 _18120_ (.A(net1248),
    .B(net818),
    .C(net1712),
    .X(_03662_));
 or2_1 _18121_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[3] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[4] ),
    .X(_03663_));
 nor2_1 _18122_ (.A(_03662_),
    .B(_03663_),
    .Y(_03664_));
 or2_1 _18123_ (.A(_03662_),
    .B(_03663_),
    .X(_03665_));
 and2_1 _18124_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[0] ),
    .B(net1176),
    .X(_03666_));
 nand2_1 _18125_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[0] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[2] ),
    .Y(_03667_));
 or2_1 _18126_ (.A(net1177),
    .B(_03667_),
    .X(_03668_));
 nor2_1 _18127_ (.A(_03665_),
    .B(_03668_),
    .Y(_03669_));
 mux2_1 _18128_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[6] ),
    .A1(net815),
    .S(_03669_),
    .X(_00468_));
 nor2_1 _18129_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[0] ),
    .B(net1176),
    .Y(_03670_));
 or3_2 _18130_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[0] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[1] ),
    .C(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[2] ),
    .X(_03671_));
 inv_2 _18131_ (.A(_03671_),
    .Y(_03672_));
 nor2_1 _18132_ (.A(_03665_),
    .B(_03671_),
    .Y(_03673_));
 mux2_1 _18133_ (.A0(\digitop_pav2.dr ),
    .A1(net816),
    .S(_03673_),
    .X(_00469_));
 and2_1 _18134_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[0] ),
    .B(_07134_),
    .X(_03674_));
 or3b_2 _18135_ (.A(net1177),
    .B(net1176),
    .C_N(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[0] ),
    .X(_03675_));
 nor2_1 _18136_ (.A(_03665_),
    .B(_03675_),
    .Y(_03676_));
 mux2_1 _18137_ (.A0(net1180),
    .A1(net816),
    .S(_03676_),
    .X(_00470_));
 and3_1 _18138_ (.A(net1177),
    .B(_03664_),
    .C(_03674_),
    .X(_03677_));
 mux2_1 _18139_ (.A0(net1179),
    .A1(net816),
    .S(_03677_),
    .X(_00471_));
 nor2_1 _18140_ (.A(_10335_),
    .B(_03665_),
    .Y(_03678_));
 mux2_1 _18141_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[3] ),
    .A1(net815),
    .S(_03678_),
    .X(_00472_));
 and3_1 _18142_ (.A(net1176),
    .B(_10334_),
    .C(_03664_),
    .X(_03679_));
 mux2_1 _18143_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[4] ),
    .A1(net816),
    .S(_03679_),
    .X(_00473_));
 and3_1 _18144_ (.A(net1177),
    .B(_03664_),
    .C(_03666_),
    .X(_03680_));
 mux2_1 _18145_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[5] ),
    .A1(net815),
    .S(_03680_),
    .X(_00474_));
 nor2_1 _18146_ (.A(_10333_),
    .B(_03662_),
    .Y(_03681_));
 or2_1 _18147_ (.A(_10333_),
    .B(_03662_),
    .X(_03682_));
 nor2_1 _18148_ (.A(_03668_),
    .B(_03682_),
    .Y(_03683_));
 mux2_1 _18149_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[1] ),
    .A1(net816),
    .S(_03683_),
    .X(_00475_));
 nor2_1 _18150_ (.A(_10333_),
    .B(_03671_),
    .Y(_03684_));
 nand2_1 _18151_ (.A(net802),
    .B(_03684_),
    .Y(_03685_));
 mux2_1 _18152_ (.A0(net815),
    .A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[7] ),
    .S(_03685_),
    .X(_00476_));
 nor2_1 _18153_ (.A(_03675_),
    .B(_03682_),
    .Y(_03686_));
 mux2_1 _18154_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[6] ),
    .A1(net814),
    .S(_03686_),
    .X(_00477_));
 and3_1 _18155_ (.A(net1177),
    .B(_03674_),
    .C(_03681_),
    .X(_03687_));
 mux2_1 _18156_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[5] ),
    .A1(net814),
    .S(_03687_),
    .X(_00478_));
 nand2_1 _18157_ (.A(_10336_),
    .B(net802),
    .Y(_03688_));
 mux2_1 _18158_ (.A0(net816),
    .A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[4] ),
    .S(_03688_),
    .X(_00479_));
 and3_1 _18159_ (.A(net1176),
    .B(_10334_),
    .C(_03681_),
    .X(_03689_));
 mux2_1 _18160_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[3] ),
    .A1(net814),
    .S(_03689_),
    .X(_00480_));
 and3_1 _18161_ (.A(net1177),
    .B(_03666_),
    .C(_03681_),
    .X(_03690_));
 mux2_1 _18162_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[2] ),
    .A1(net815),
    .S(_03690_),
    .X(_00481_));
 nor2_1 _18163_ (.A(_10340_),
    .B(_03662_),
    .Y(_03691_));
 or2_1 _18164_ (.A(_10340_),
    .B(_03662_),
    .X(_03692_));
 nor2_1 _18165_ (.A(_03668_),
    .B(_03692_),
    .Y(_03693_));
 mux2_1 _18166_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[6] ),
    .A1(net814),
    .S(_03693_),
    .X(_00482_));
 nor2_1 _18167_ (.A(_03671_),
    .B(_03692_),
    .Y(_03694_));
 mux2_1 _18168_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[0] ),
    .A1(net815),
    .S(_03694_),
    .X(_00483_));
 nor2_1 _18169_ (.A(_03675_),
    .B(_03692_),
    .Y(_03695_));
 mux2_1 _18170_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[1] ),
    .A1(net814),
    .S(_03695_),
    .X(_00484_));
 and3_1 _18171_ (.A(net1177),
    .B(_03674_),
    .C(_03691_),
    .X(_03696_));
 mux2_1 _18172_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[2] ),
    .A1(net815),
    .S(_03696_),
    .X(_00485_));
 nor2_1 _18173_ (.A(_10335_),
    .B(_03692_),
    .Y(_03697_));
 mux2_1 _18174_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[3] ),
    .A1(net814),
    .S(_03697_),
    .X(_00486_));
 and3_1 _18175_ (.A(net1176),
    .B(_10334_),
    .C(_03691_),
    .X(_03698_));
 mux2_1 _18176_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[4] ),
    .A1(net814),
    .S(_03698_),
    .X(_00487_));
 and3_1 _18177_ (.A(net1177),
    .B(_03666_),
    .C(_03691_),
    .X(_03699_));
 mux2_1 _18178_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[5] ),
    .A1(net814),
    .S(_03699_),
    .X(_00488_));
 o21ba_1 _18179_ (.A1(s1_set_ff2),
    .A2(\digitop_pav2.s1_i ),
    .B1_N(net1837),
    .X(_00489_));
 or4b_4 _18180_ (.A(\digitop_pav2.sec_inst.shift_in.st[0] ),
    .B(\digitop_pav2.sec_inst.shift_in.st[1] ),
    .C(_11400_),
    .D_N(\digitop_pav2.sec_inst.shift_in.st[4] ),
    .X(_03700_));
 o21ba_1 _18181_ (.A1(net717),
    .A2(\digitop_pav2.sec_inst.ld_r.st[0] ),
    .B1_N(\digitop_pav2.sec_inst.ld_r.st[1] ),
    .X(_03701_));
 a2111o_1 _18182_ (.A1(\digitop_pav2.sec_inst.sm.st[6] ),
    .A2(net366),
    .B1(_09652_),
    .C1(_03700_),
    .D1(_03701_),
    .X(_03702_));
 a211o_1 _18183_ (.A1(net1652),
    .A2(\digitop_pav2.sec_inst.sm.st[1] ),
    .B1(_03702_),
    .C1(\digitop_pav2.sec_inst.en_shifto ),
    .X(_03703_));
 inv_2 _18184_ (.A(_03703_),
    .Y(_03704_));
 a21oi_4 _18185_ (.A1(\digitop_pav2.sec_inst.sm.st[9] ),
    .A2(net1646),
    .B1(_03703_),
    .Y(_03705_));
 a21o_2 _18186_ (.A1(\digitop_pav2.sec_inst.sm.st[9] ),
    .A2(net1646),
    .B1(_03703_),
    .X(_03706_));
 and2_1 _18187_ (.A(\digitop_pav2.sec_inst.sm.next_st[1] ),
    .B(net1647),
    .X(_00490_));
 mux2_1 _18188_ (.A0(\digitop_pav2.sec_inst.sm.st[1] ),
    .A1(\digitop_pav2.sec_inst.sm.next_st[1] ),
    .S(net1653),
    .X(_00491_));
 a311o_1 _18189_ (.A1(\digitop_pav2.sec_inst.en_ld_data ),
    .A2(net702),
    .A3(_07107_),
    .B1(\digitop_pav2.sec_inst.sm.st[1] ),
    .C1(net719),
    .X(_03707_));
 and3b_1 _18190_ (.A_N(\digitop_pav2.sec_inst.sm.st[1] ),
    .B(net1621),
    .C(net719),
    .X(_03708_));
 or4b_1 _18191_ (.A(\digitop_pav2.sec_inst.sm.next_st[1] ),
    .B(_03708_),
    .C(net1647),
    .D_N(_03707_),
    .X(_03709_));
 a21bo_1 _18192_ (.A1(net719),
    .A2(net1647),
    .B1_N(_03709_),
    .X(_00492_));
 and3b_1 _18193_ (.A_N(\digitop_pav2.sec_inst.sm.next_st[1] ),
    .B(net1653),
    .C(_03708_),
    .X(_03710_));
 a21o_1 _18194_ (.A1(\digitop_pav2.rng_inst.rng_prngx_pav2.rngx_sec_req_i ),
    .A2(net1647),
    .B1(_03710_),
    .X(_00493_));
 nor2_1 _18195_ (.A(\digitop_pav2.sec_inst.sm.st[6] ),
    .B(_09166_),
    .Y(_03711_));
 and3b_1 _18196_ (.A_N(\digitop_pav2.sec_inst.sm.st[9] ),
    .B(net712),
    .C(_03711_),
    .X(_03712_));
 a311o_1 _18197_ (.A1(net715),
    .A2(_07064_),
    .A3(_03702_),
    .B1(_03712_),
    .C1(\digitop_pav2.rng_inst.rng_prngx_pav2.rngx_sec_req_i ),
    .X(_03713_));
 or3_1 _18198_ (.A(net719),
    .B(\digitop_pav2.sec_inst.sm.st[1] ),
    .C(\digitop_pav2.sec_inst.sm.next_st[1] ),
    .X(_03714_));
 nand2_1 _18199_ (.A(_07064_),
    .B(net1006),
    .Y(_03715_));
 nor2_1 _18200_ (.A(\digitop_pav2.rng_inst.rng_prngx_pav2.rngx_sec_req_i ),
    .B(_03714_),
    .Y(_03716_));
 nor2_1 _18201_ (.A(_03714_),
    .B(_03715_),
    .Y(_03717_));
 o21a_1 _18202_ (.A1(_03716_),
    .A2(_03717_),
    .B1(_03713_),
    .X(_03718_));
 mux2_1 _18203_ (.A0(net715),
    .A1(_03718_),
    .S(net1653),
    .X(_00494_));
 or4b_1 _18204_ (.A(net702),
    .B(\digitop_pav2.rng_inst.rng_prngx_pav2.rngx_sec_req_i ),
    .C(_03702_),
    .D_N(net715),
    .X(_03719_));
 or3_1 _18205_ (.A(_07064_),
    .B(_07107_),
    .C(net1624),
    .X(_03720_));
 a21o_1 _18206_ (.A1(_03719_),
    .A2(_03720_),
    .B1(net1647),
    .X(_03721_));
 a2bb2o_1 _18207_ (.A1_N(_03714_),
    .A2_N(_03721_),
    .B1(\digitop_pav2.sec_inst.dg_key.en_i ),
    .B2(net1647),
    .X(_00495_));
 nand2_1 _18208_ (.A(net1653),
    .B(_03716_),
    .Y(_03722_));
 a2bb2o_1 _18209_ (.A1_N(_09655_),
    .A2_N(_03722_),
    .B1(net1647),
    .B2(\digitop_pav2.sec_inst.sm.st[6] ),
    .X(_00496_));
 a41o_1 _18210_ (.A1(\digitop_pav2.sec_inst.sm.st[9] ),
    .A2(net1653),
    .A3(_03711_),
    .A4(_03716_),
    .B1(\digitop_pav2.sec_inst.en_shifto ),
    .X(_00497_));
 nand2_1 _18211_ (.A(\digitop_pav2.sec_inst.sm.st[6] ),
    .B(_03716_),
    .Y(_03723_));
 or4_1 _18212_ (.A(_09166_),
    .B(net1647),
    .C(_03715_),
    .D(_03723_),
    .X(_03724_));
 o21ai_1 _18213_ (.A1(net697),
    .A2(net1653),
    .B1(_03724_),
    .Y(_00498_));
 a41o_1 _18214_ (.A1(\digitop_pav2.sec_inst.sm.st[6] ),
    .A2(_09165_),
    .A3(_03715_),
    .A4(_03716_),
    .B1(net1647),
    .X(_03725_));
 o21a_1 _18215_ (.A1(\digitop_pav2.sec_inst.sm.st[9] ),
    .A2(_03704_),
    .B1(_03725_),
    .X(_00499_));
 and2_1 _18216_ (.A(net1446),
    .B(\digitop_pav2.sync_inst.inst_rstx.gray_counter[1] ),
    .X(_03726_));
 a31o_1 _18217_ (.A1(net1400),
    .A2(_07236_),
    .A3(\digitop_pav2.sync_inst.inst_rstx.gray_counter[0] ),
    .B1(_03726_),
    .X(_00500_));
 a21o_1 _18218_ (.A1(net1400),
    .A2(\digitop_pav2.sync_inst.inst_rstx.gray_counter[1] ),
    .B1(\digitop_pav2.sync_inst.inst_rstx.gray_counter[2] ),
    .X(_03727_));
 o21a_1 _18219_ (.A1(net1446),
    .A2(\digitop_pav2.sync_inst.inst_rstx.gray_counter[0] ),
    .B1(_03727_),
    .X(_00501_));
 a211o_1 _18220_ (.A1(_07055_),
    .A2(_07156_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[2] ),
    .C1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[4] ),
    .X(_03728_));
 a21oi_1 _18221_ (.A1(_07055_),
    .A2(_09635_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_read ),
    .Y(_03729_));
 and2_1 _18222_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[0] ),
    .B(_03729_),
    .X(_03730_));
 nor3_1 _18223_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[4] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[2] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[3] ),
    .Y(_03731_));
 nand2_1 _18224_ (.A(_07055_),
    .B(net1473),
    .Y(_03732_));
 inv_2 _18225_ (.A(_03732_),
    .Y(_03733_));
 a21o_1 _18226_ (.A1(_09634_),
    .A2(_09636_),
    .B1(_03732_),
    .X(_03734_));
 mux2_1 _18227_ (.A0(_09631_),
    .A1(net1473),
    .S(_07055_),
    .X(_03735_));
 a211o_1 _18228_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[2] ),
    .A2(_09634_),
    .B1(_09641_),
    .C1(_03735_),
    .X(_03736_));
 nand2_2 _18229_ (.A(_03734_),
    .B(_03736_),
    .Y(_03737_));
 or2_1 _18230_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[0] ),
    .B(_03729_),
    .X(_03738_));
 nand2_1 _18231_ (.A(_03737_),
    .B(_03738_),
    .Y(_03739_));
 o32a_1 _18232_ (.A1(_09629_),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_read ),
    .A3(_03728_),
    .B1(_03730_),
    .B2(_03739_),
    .X(_00502_));
 o21ai_1 _18233_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[1] ),
    .A2(_03738_),
    .B1(_03737_),
    .Y(_03740_));
 a21o_1 _18234_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[1] ),
    .A2(_03738_),
    .B1(_03740_),
    .X(_00503_));
 o31a_1 _18235_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[1] ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[2] ),
    .A3(_03738_),
    .B1(_03737_),
    .X(_03741_));
 a21o_1 _18236_ (.A1(_09640_),
    .A2(_03731_),
    .B1(_03741_),
    .X(_03742_));
 o21ai_1 _18237_ (.A1(_07154_),
    .A2(_03740_),
    .B1(_03742_),
    .Y(_00504_));
 a21o_1 _18238_ (.A1(_03729_),
    .A2(_03737_),
    .B1(_09632_),
    .X(_03743_));
 a211o_1 _18239_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[2] ),
    .A2(_09635_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_read ),
    .C1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[4] ),
    .X(_03744_));
 or3_1 _18240_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[0] ),
    .B(net1473),
    .C(_03744_),
    .X(_03745_));
 or3_1 _18241_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[3] ),
    .B(_09632_),
    .C(_03729_),
    .X(_03746_));
 nand2_1 _18242_ (.A(_03737_),
    .B(_03746_),
    .Y(_03747_));
 a22o_1 _18243_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[3] ),
    .A2(_03743_),
    .B1(_03745_),
    .B2(_03747_),
    .X(_00505_));
 and2_1 _18244_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[4] ),
    .B(_03746_),
    .X(_03748_));
 o21ai_1 _18245_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[4] ),
    .A2(_03746_),
    .B1(_03737_),
    .Y(_03749_));
 o32a_1 _18246_ (.A1(_09629_),
    .A2(_03733_),
    .A3(_03744_),
    .B1(_03748_),
    .B2(_03749_),
    .X(_00506_));
 a21bo_1 _18247_ (.A1(_09634_),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_read ),
    .B1_N(_03737_),
    .X(_03750_));
 a211o_1 _18248_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[0] ),
    .A2(_09630_),
    .B1(_03737_),
    .C1(_03744_),
    .X(_03751_));
 a2bb2o_1 _18249_ (.A1_N(_07155_),
    .A2_N(_03749_),
    .B1(_03750_),
    .B2(_03751_),
    .X(_00507_));
 nand2_1 _18250_ (.A(_09634_),
    .B(_03733_),
    .Y(_03752_));
 a21oi_2 _18251_ (.A1(_09634_),
    .A2(_03733_),
    .B1(_09628_),
    .Y(_03753_));
 o21ai_2 _18252_ (.A1(_07156_),
    .A2(_11108_),
    .B1(_03753_),
    .Y(_03754_));
 o21ai_2 _18253_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.int_wr_bit ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_bit ),
    .B1(_09628_),
    .Y(_03755_));
 nand2_1 _18254_ (.A(net1460),
    .B(_03755_),
    .Y(_03756_));
 and2_1 _18255_ (.A(net1478),
    .B(net1477),
    .X(_03757_));
 nand2_1 _18256_ (.A(net1478),
    .B(net1477),
    .Y(_03758_));
 a22o_4 _18257_ (.A1(_09403_),
    .A2(_09405_),
    .B1(_09416_),
    .B2(net957),
    .X(_03759_));
 o2bb2a_2 _18258_ (.A1_N(_09403_),
    .A2_N(_09405_),
    .B1(_09415_),
    .B2(_09388_),
    .X(_03760_));
 or2_1 _18259_ (.A(_09387_),
    .B(_09391_),
    .X(_03761_));
 nor2_1 _18260_ (.A(_09387_),
    .B(_09391_),
    .Y(_03762_));
 mux2_1 _18261_ (.A0(\vmem_after_buf[320] ),
    .A1(\vmem_after_buf[336] ),
    .S(net952),
    .X(_03763_));
 or4_1 _18262_ (.A(net120),
    .B(net121),
    .C(net122),
    .D(net123),
    .X(_03764_));
 nor4_1 _18263_ (.A(_11005_),
    .B(_11007_),
    .C(_11010_),
    .D(_03764_),
    .Y(_03765_));
 or4_4 _18264_ (.A(_11005_),
    .B(_11007_),
    .C(_11010_),
    .D(_03764_),
    .X(_03766_));
 mux2_1 _18265_ (.A0(\vmem_after_buf[352] ),
    .A1(\vmem_after_buf[368] ),
    .S(net952),
    .X(_03767_));
 mux2_1 _18266_ (.A0(_03763_),
    .A1(_03767_),
    .S(net891),
    .X(_03768_));
 mux2_1 _18267_ (.A0(\vmem_after_buf[256] ),
    .A1(\vmem_after_buf[272] ),
    .S(net952),
    .X(_03769_));
 mux2_1 _18268_ (.A0(\vmem_after_buf[288] ),
    .A1(\vmem_after_buf[304] ),
    .S(net952),
    .X(_03770_));
 mux2_1 _18269_ (.A0(_03769_),
    .A1(_03770_),
    .S(net891),
    .X(_03771_));
 mux2_1 _18270_ (.A0(_03768_),
    .A1(_03771_),
    .S(net767),
    .X(_03772_));
 mux2_1 _18271_ (.A0(net27),
    .A1(_03772_),
    .S(net1493),
    .X(_03773_));
 mux2_1 _18272_ (.A0(\vmem_after_buf[80] ),
    .A1(\vmem_after_buf[64] ),
    .S(net923),
    .X(_03774_));
 mux2_1 _18273_ (.A0(\vmem_after_buf[112] ),
    .A1(\vmem_after_buf[96] ),
    .S(net923),
    .X(_03775_));
 mux2_1 _18274_ (.A0(_03774_),
    .A1(_03775_),
    .S(net891),
    .X(_03776_));
 mux2_1 _18275_ (.A0(\vmem_after_buf[16] ),
    .A1(\vmem_after_buf[0] ),
    .S(net923),
    .X(_03777_));
 mux2_1 _18276_ (.A0(\vmem_after_buf[48] ),
    .A1(\vmem_after_buf[32] ),
    .S(net923),
    .X(_03778_));
 mux2_1 _18277_ (.A0(_03777_),
    .A1(_03778_),
    .S(net891),
    .X(_03779_));
 mux2_1 _18278_ (.A0(_03776_),
    .A1(_03779_),
    .S(net766),
    .X(_03780_));
 mux2_1 _18279_ (.A0(net2),
    .A1(_03780_),
    .S(net1493),
    .X(_03781_));
 nor2_1 _18280_ (.A(net1478),
    .B(net1477),
    .Y(_03782_));
 mux2_1 _18281_ (.A0(\vmem_after_buf[208] ),
    .A1(\vmem_after_buf[192] ),
    .S(net919),
    .X(_03783_));
 mux2_1 _18282_ (.A0(\vmem_after_buf[240] ),
    .A1(\vmem_after_buf[224] ),
    .S(net919),
    .X(_03784_));
 mux2_1 _18283_ (.A0(_03783_),
    .A1(_03784_),
    .S(net889),
    .X(_03785_));
 mux2_1 _18284_ (.A0(\vmem_after_buf[144] ),
    .A1(\vmem_after_buf[128] ),
    .S(net919),
    .X(_03786_));
 mux2_1 _18285_ (.A0(\vmem_after_buf[176] ),
    .A1(\vmem_after_buf[160] ),
    .S(net919),
    .X(_03787_));
 mux2_1 _18286_ (.A0(_03786_),
    .A1(_03787_),
    .S(net889),
    .X(_03788_));
 mux2_1 _18287_ (.A0(_03785_),
    .A1(_03788_),
    .S(net762),
    .X(_03789_));
 mux2_1 _18288_ (.A0(net9),
    .A1(_03789_),
    .S(net1493),
    .X(_03790_));
 a22o_1 _18289_ (.A1(net1477),
    .A2(_03773_),
    .B1(_03790_),
    .B2(net1478),
    .X(_03791_));
 a211o_1 _18290_ (.A1(_03781_),
    .A2(net1468),
    .B1(_03791_),
    .C1(net1472),
    .X(_03792_));
 mux2_1 _18291_ (.A0(\vmem_after_buf[448] ),
    .A1(\vmem_after_buf[464] ),
    .S(net955),
    .X(_03793_));
 mux2_1 _18292_ (.A0(\vmem_after_buf[480] ),
    .A1(\vmem_after_buf[496] ),
    .S(net952),
    .X(_03794_));
 mux2_1 _18293_ (.A0(_03793_),
    .A1(_03794_),
    .S(net891),
    .X(_03795_));
 mux2_1 _18294_ (.A0(\vmem_after_buf[384] ),
    .A1(\vmem_after_buf[400] ),
    .S(net955),
    .X(_03796_));
 mux2_1 _18295_ (.A0(\vmem_after_buf[416] ),
    .A1(\vmem_after_buf[432] ),
    .S(net952),
    .X(_03797_));
 mux2_1 _18296_ (.A0(_03796_),
    .A1(_03797_),
    .S(net891),
    .X(_03798_));
 mux2_1 _18297_ (.A0(_03795_),
    .A1(_03798_),
    .S(net767),
    .X(_03799_));
 mux2_1 _18298_ (.A0(net44),
    .A1(_03799_),
    .S(net1493),
    .X(_03800_));
 o211a_1 _18299_ (.A1(_03758_),
    .A2(_03800_),
    .B1(_03792_),
    .C1(net1463),
    .X(_03801_));
 o22a_1 _18300_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[0] ),
    .A2(net1460),
    .B1(net1394),
    .B2(_03801_),
    .X(_00508_));
 mux2_1 _18301_ (.A0(\vmem_after_buf[49] ),
    .A1(\vmem_after_buf[33] ),
    .S(net939),
    .X(_03802_));
 mux2_1 _18302_ (.A0(\vmem_after_buf[17] ),
    .A1(\vmem_after_buf[1] ),
    .S(net940),
    .X(_03803_));
 mux2_1 _18303_ (.A0(_03802_),
    .A1(_03803_),
    .S(net910),
    .X(_03804_));
 mux2_1 _18304_ (.A0(\vmem_after_buf[81] ),
    .A1(\vmem_after_buf[65] ),
    .S(net941),
    .X(_03805_));
 mux2_1 _18305_ (.A0(\vmem_after_buf[113] ),
    .A1(\vmem_after_buf[97] ),
    .S(net943),
    .X(_03806_));
 mux2_1 _18306_ (.A0(_03805_),
    .A1(_03806_),
    .S(net900),
    .X(_03807_));
 mux2_1 _18307_ (.A0(_03804_),
    .A1(_03807_),
    .S(net743),
    .X(_03808_));
 mux2_1 _18308_ (.A0(net13),
    .A1(_03808_),
    .S(net1492),
    .X(_03809_));
 mux2_1 _18309_ (.A0(\vmem_after_buf[209] ),
    .A1(\vmem_after_buf[193] ),
    .S(net943),
    .X(_03810_));
 mux2_1 _18310_ (.A0(\vmem_after_buf[241] ),
    .A1(\vmem_after_buf[225] ),
    .S(net943),
    .X(_03811_));
 mux2_1 _18311_ (.A0(_03810_),
    .A1(_03811_),
    .S(net901),
    .X(_03812_));
 mux2_1 _18312_ (.A0(\vmem_after_buf[145] ),
    .A1(\vmem_after_buf[129] ),
    .S(net943),
    .X(_03813_));
 mux2_1 _18313_ (.A0(\vmem_after_buf[177] ),
    .A1(\vmem_after_buf[161] ),
    .S(net943),
    .X(_03814_));
 mux2_1 _18314_ (.A0(_03813_),
    .A1(_03814_),
    .S(net901),
    .X(_03815_));
 mux2_1 _18315_ (.A0(_03812_),
    .A1(_03815_),
    .S(net791),
    .X(_03816_));
 mux2_1 _18316_ (.A0(net10),
    .A1(_03816_),
    .S(net1492),
    .X(_03817_));
 mux2_1 _18317_ (.A0(\vmem_after_buf[337] ),
    .A1(\vmem_after_buf[321] ),
    .S(net942),
    .X(_03818_));
 mux2_1 _18318_ (.A0(\vmem_after_buf[369] ),
    .A1(\vmem_after_buf[353] ),
    .S(net942),
    .X(_03819_));
 mux2_1 _18319_ (.A0(_03818_),
    .A1(_03819_),
    .S(net905),
    .X(_03820_));
 mux2_1 _18320_ (.A0(\vmem_after_buf[273] ),
    .A1(\vmem_after_buf[257] ),
    .S(net942),
    .X(_03821_));
 mux2_1 _18321_ (.A0(\vmem_after_buf[305] ),
    .A1(\vmem_after_buf[289] ),
    .S(net942),
    .X(_03822_));
 mux2_1 _18322_ (.A0(_03821_),
    .A1(_03822_),
    .S(net901),
    .X(_03823_));
 mux2_1 _18323_ (.A0(_03820_),
    .A1(_03823_),
    .S(net789),
    .X(_03824_));
 mux2_1 _18324_ (.A0(net28),
    .A1(_03824_),
    .S(net1493),
    .X(_03825_));
 and2b_1 _18325_ (.A_N(net1478),
    .B(net1477),
    .X(_03826_));
 a22o_1 _18326_ (.A1(net1469),
    .A2(_03809_),
    .B1(_03825_),
    .B2(net1467),
    .X(_03827_));
 and2b_2 _18327_ (.A_N(net1477),
    .B(net1478),
    .X(_03828_));
 a211o_1 _18328_ (.A1(net1478),
    .A2(_03817_),
    .B1(_03827_),
    .C1(net1471),
    .X(_03829_));
 mux2_1 _18329_ (.A0(\vmem_after_buf[433] ),
    .A1(\vmem_after_buf[417] ),
    .S(net943),
    .X(_03830_));
 mux2_1 _18330_ (.A0(\vmem_after_buf[401] ),
    .A1(\vmem_after_buf[385] ),
    .S(net942),
    .X(_03831_));
 mux2_1 _18331_ (.A0(_03830_),
    .A1(_03831_),
    .S(net910),
    .X(_03832_));
 mux2_1 _18332_ (.A0(\vmem_after_buf[465] ),
    .A1(\vmem_after_buf[449] ),
    .S(net942),
    .X(_03833_));
 mux2_1 _18333_ (.A0(\vmem_after_buf[497] ),
    .A1(\vmem_after_buf[481] ),
    .S(net943),
    .X(_03834_));
 mux2_1 _18334_ (.A0(_03833_),
    .A1(_03834_),
    .S(net901),
    .X(_03835_));
 mux2_1 _18335_ (.A0(_03832_),
    .A1(_03835_),
    .S(net746),
    .X(_03836_));
 mux2_2 _18336_ (.A0(net45),
    .A1(_03836_),
    .S(net1499),
    .X(_03837_));
 o211a_1 _18337_ (.A1(_03758_),
    .A2(_03837_),
    .B1(_03829_),
    .C1(net1462),
    .X(_03838_));
 nor2_1 _18338_ (.A(_09628_),
    .B(_03752_),
    .Y(_03839_));
 a21o_1 _18339_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[0] ),
    .A2(net1458),
    .B1(net1395),
    .X(_03840_));
 o22a_1 _18340_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[1] ),
    .A2(net1461),
    .B1(_03838_),
    .B2(_03840_),
    .X(_00509_));
 mux2_1 _18341_ (.A0(\vmem_after_buf[82] ),
    .A1(\vmem_after_buf[66] ),
    .S(net944),
    .X(_03841_));
 mux2_1 _18342_ (.A0(\vmem_after_buf[114] ),
    .A1(\vmem_after_buf[98] ),
    .S(net944),
    .X(_03842_));
 mux2_1 _18343_ (.A0(_03841_),
    .A1(_03842_),
    .S(net902),
    .X(_03843_));
 mux2_1 _18344_ (.A0(\vmem_after_buf[18] ),
    .A1(\vmem_after_buf[2] ),
    .S(net944),
    .X(_03844_));
 mux2_1 _18345_ (.A0(\vmem_after_buf[50] ),
    .A1(\vmem_after_buf[34] ),
    .S(net944),
    .X(_03845_));
 mux2_1 _18346_ (.A0(_03844_),
    .A1(_03845_),
    .S(net902),
    .X(_03846_));
 mux2_1 _18347_ (.A0(_03843_),
    .A1(_03846_),
    .S(net792),
    .X(_03847_));
 mux2_1 _18348_ (.A0(net24),
    .A1(_03847_),
    .S(net1498),
    .X(_03848_));
 mux2_1 _18349_ (.A0(\vmem_after_buf[338] ),
    .A1(\vmem_after_buf[322] ),
    .S(net940),
    .X(_03849_));
 mux2_1 _18350_ (.A0(\vmem_after_buf[370] ),
    .A1(\vmem_after_buf[354] ),
    .S(net941),
    .X(_03850_));
 mux2_1 _18351_ (.A0(_03849_),
    .A1(_03850_),
    .S(net900),
    .X(_03851_));
 mux2_1 _18352_ (.A0(\vmem_after_buf[274] ),
    .A1(\vmem_after_buf[258] ),
    .S(net940),
    .X(_03852_));
 mux2_1 _18353_ (.A0(\vmem_after_buf[306] ),
    .A1(\vmem_after_buf[290] ),
    .S(net940),
    .X(_03853_));
 mux2_1 _18354_ (.A0(_03852_),
    .A1(_03853_),
    .S(net901),
    .X(_03854_));
 mux2_1 _18355_ (.A0(_03851_),
    .A1(_03854_),
    .S(net787),
    .X(_03855_));
 mux2_1 _18356_ (.A0(net29),
    .A1(_03855_),
    .S(net1495),
    .X(_03856_));
 mux2_1 _18357_ (.A0(\vmem_after_buf[178] ),
    .A1(\vmem_after_buf[162] ),
    .S(net940),
    .X(_03857_));
 mux2_1 _18358_ (.A0(\vmem_after_buf[146] ),
    .A1(\vmem_after_buf[130] ),
    .S(net940),
    .X(_03858_));
 mux2_1 _18359_ (.A0(_03857_),
    .A1(_03858_),
    .S(net910),
    .X(_03859_));
 mux2_1 _18360_ (.A0(\vmem_after_buf[210] ),
    .A1(\vmem_after_buf[194] ),
    .S(net940),
    .X(_03860_));
 mux2_1 _18361_ (.A0(\vmem_after_buf[242] ),
    .A1(\vmem_after_buf[226] ),
    .S(net940),
    .X(_03861_));
 mux2_1 _18362_ (.A0(_03860_),
    .A1(_03861_),
    .S(net901),
    .X(_03862_));
 mux2_1 _18363_ (.A0(_03859_),
    .A1(_03862_),
    .S(net745),
    .X(_03863_));
 mux2_1 _18364_ (.A0(net11),
    .A1(_03863_),
    .S(net1496),
    .X(_03864_));
 a22o_1 _18365_ (.A1(net1469),
    .A2(_03848_),
    .B1(_03856_),
    .B2(net1477),
    .X(_03865_));
 a211o_1 _18366_ (.A1(net1478),
    .A2(_03864_),
    .B1(_03865_),
    .C1(net1471),
    .X(_03866_));
 mux2_1 _18367_ (.A0(\vmem_after_buf[466] ),
    .A1(\vmem_after_buf[450] ),
    .S(net944),
    .X(_03867_));
 mux2_1 _18368_ (.A0(\vmem_after_buf[498] ),
    .A1(\vmem_after_buf[482] ),
    .S(net946),
    .X(_03868_));
 mux2_1 _18369_ (.A0(_03867_),
    .A1(_03868_),
    .S(net902),
    .X(_03869_));
 mux2_1 _18370_ (.A0(\vmem_after_buf[402] ),
    .A1(\vmem_after_buf[386] ),
    .S(net944),
    .X(_03870_));
 mux2_1 _18371_ (.A0(\vmem_after_buf[434] ),
    .A1(\vmem_after_buf[418] ),
    .S(net944),
    .X(_03871_));
 mux2_1 _18372_ (.A0(_03870_),
    .A1(_03871_),
    .S(net902),
    .X(_03872_));
 mux2_1 _18373_ (.A0(_03869_),
    .A1(_03872_),
    .S(net795),
    .X(_03873_));
 mux2_1 _18374_ (.A0(net47),
    .A1(_03873_),
    .S(net1499),
    .X(_03874_));
 o211a_1 _18375_ (.A1(net1470),
    .A2(_03874_),
    .B1(_03866_),
    .C1(net1462),
    .X(_03875_));
 a21o_1 _18376_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[1] ),
    .A2(net1459),
    .B1(net1395),
    .X(_03876_));
 o22a_1 _18377_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[2] ),
    .A2(net1461),
    .B1(_03875_),
    .B2(_03876_),
    .X(_00510_));
 mux2_1 _18378_ (.A0(\vmem_after_buf[51] ),
    .A1(\vmem_after_buf[35] ),
    .S(net918),
    .X(_03877_));
 mux2_1 _18379_ (.A0(\vmem_after_buf[19] ),
    .A1(\vmem_after_buf[3] ),
    .S(net916),
    .X(_03878_));
 mux2_1 _18380_ (.A0(_03877_),
    .A1(_03878_),
    .S(net906),
    .X(_03879_));
 mux2_1 _18381_ (.A0(\vmem_after_buf[83] ),
    .A1(\vmem_after_buf[67] ),
    .S(net918),
    .X(_03880_));
 mux2_1 _18382_ (.A0(\vmem_after_buf[115] ),
    .A1(\vmem_after_buf[99] ),
    .S(net916),
    .X(_03881_));
 mux2_1 _18383_ (.A0(_03880_),
    .A1(_03881_),
    .S(net887),
    .X(_03882_));
 mux2_1 _18384_ (.A0(_03879_),
    .A1(_03882_),
    .S(net722),
    .X(_03883_));
 mux2_1 _18385_ (.A0(net35),
    .A1(_03883_),
    .S(net1494),
    .X(_03884_));
 mux2_1 _18386_ (.A0(\vmem_after_buf[211] ),
    .A1(\vmem_after_buf[195] ),
    .S(net916),
    .X(_03885_));
 mux2_1 _18387_ (.A0(\vmem_after_buf[243] ),
    .A1(\vmem_after_buf[227] ),
    .S(net916),
    .X(_03886_));
 mux2_1 _18388_ (.A0(_03885_),
    .A1(_03886_),
    .S(net887),
    .X(_03887_));
 mux2_1 _18389_ (.A0(\vmem_after_buf[147] ),
    .A1(\vmem_after_buf[131] ),
    .S(net916),
    .X(_03888_));
 mux2_1 _18390_ (.A0(\vmem_after_buf[179] ),
    .A1(\vmem_after_buf[163] ),
    .S(net916),
    .X(_03889_));
 mux2_1 _18391_ (.A0(_03888_),
    .A1(_03889_),
    .S(net887),
    .X(_03890_));
 mux2_1 _18392_ (.A0(_03887_),
    .A1(_03890_),
    .S(net758),
    .X(_03891_));
 mux2_1 _18393_ (.A0(net12),
    .A1(_03891_),
    .S(net1494),
    .X(_03892_));
 mux2_1 _18394_ (.A0(\vmem_after_buf[339] ),
    .A1(\vmem_after_buf[323] ),
    .S(net917),
    .X(_03893_));
 mux2_1 _18395_ (.A0(\vmem_after_buf[371] ),
    .A1(\vmem_after_buf[355] ),
    .S(net916),
    .X(_03894_));
 mux2_1 _18396_ (.A0(_03893_),
    .A1(_03894_),
    .S(net888),
    .X(_03895_));
 mux2_1 _18397_ (.A0(\vmem_after_buf[275] ),
    .A1(\vmem_after_buf[259] ),
    .S(net917),
    .X(_03896_));
 mux2_1 _18398_ (.A0(\vmem_after_buf[307] ),
    .A1(\vmem_after_buf[291] ),
    .S(net917),
    .X(_03897_));
 mux2_1 _18399_ (.A0(_03896_),
    .A1(_03897_),
    .S(net888),
    .X(_03898_));
 mux2_1 _18400_ (.A0(_03895_),
    .A1(_03898_),
    .S(net760),
    .X(_03899_));
 mux2_1 _18401_ (.A0(net30),
    .A1(_03899_),
    .S(net1492),
    .X(_03900_));
 a22o_1 _18402_ (.A1(_03828_),
    .A2(_03892_),
    .B1(_03900_),
    .B2(net1467),
    .X(_03901_));
 a211o_1 _18403_ (.A1(net1468),
    .A2(_03884_),
    .B1(_03901_),
    .C1(net1472),
    .X(_03902_));
 mux2_1 _18404_ (.A0(\vmem_after_buf[467] ),
    .A1(\vmem_after_buf[451] ),
    .S(net916),
    .X(_03903_));
 mux2_1 _18405_ (.A0(\vmem_after_buf[499] ),
    .A1(\vmem_after_buf[483] ),
    .S(net916),
    .X(_03904_));
 mux2_1 _18406_ (.A0(_03903_),
    .A1(_03904_),
    .S(net887),
    .X(_03905_));
 mux2_1 _18407_ (.A0(\vmem_after_buf[403] ),
    .A1(\vmem_after_buf[387] ),
    .S(net917),
    .X(_03906_));
 mux2_1 _18408_ (.A0(\vmem_after_buf[435] ),
    .A1(\vmem_after_buf[419] ),
    .S(net917),
    .X(_03907_));
 mux2_1 _18409_ (.A0(_03906_),
    .A1(_03907_),
    .S(net888),
    .X(_03908_));
 mux2_1 _18410_ (.A0(_03905_),
    .A1(_03908_),
    .S(net760),
    .X(_03909_));
 mux2_1 _18411_ (.A0(net48),
    .A1(_03909_),
    .S(net1494),
    .X(_03910_));
 o211a_1 _18412_ (.A1(net1470),
    .A2(_03910_),
    .B1(_03902_),
    .C1(net1463),
    .X(_03911_));
 a21o_1 _18413_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[2] ),
    .A2(net1458),
    .B1(net1394),
    .X(_03912_));
 o22a_1 _18414_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[3] ),
    .A2(net1460),
    .B1(_03911_),
    .B2(_03912_),
    .X(_00511_));
 mux2_1 _18415_ (.A0(\vmem_after_buf[84] ),
    .A1(\vmem_after_buf[68] ),
    .S(net945),
    .X(_03913_));
 mux2_1 _18416_ (.A0(\vmem_after_buf[116] ),
    .A1(\vmem_after_buf[100] ),
    .S(net945),
    .X(_03914_));
 mux2_1 _18417_ (.A0(_03913_),
    .A1(_03914_),
    .S(net902),
    .X(_03915_));
 mux2_1 _18418_ (.A0(\vmem_after_buf[20] ),
    .A1(\vmem_after_buf[4] ),
    .S(net945),
    .X(_03916_));
 mux2_1 _18419_ (.A0(\vmem_after_buf[52] ),
    .A1(\vmem_after_buf[36] ),
    .S(net946),
    .X(_03917_));
 mux2_1 _18420_ (.A0(_03916_),
    .A1(_03917_),
    .S(net902),
    .X(_03918_));
 mux2_1 _18421_ (.A0(_03915_),
    .A1(_03918_),
    .S(net794),
    .X(_03919_));
 mux2_2 _18422_ (.A0(net46),
    .A1(_03919_),
    .S(net1499),
    .X(_03920_));
 mux2_1 _18423_ (.A0(\vmem_after_buf[212] ),
    .A1(\vmem_after_buf[196] ),
    .S(net945),
    .X(_03921_));
 mux2_1 _18424_ (.A0(\vmem_after_buf[244] ),
    .A1(\vmem_after_buf[228] ),
    .S(net945),
    .X(_03922_));
 mux2_1 _18425_ (.A0(_03921_),
    .A1(_03922_),
    .S(net904),
    .X(_03923_));
 mux2_1 _18426_ (.A0(\vmem_after_buf[148] ),
    .A1(\vmem_after_buf[132] ),
    .S(net945),
    .X(_03924_));
 mux2_1 _18427_ (.A0(\vmem_after_buf[180] ),
    .A1(\vmem_after_buf[164] ),
    .S(net945),
    .X(_03925_));
 mux2_1 _18428_ (.A0(_03924_),
    .A1(_03925_),
    .S(net904),
    .X(_03926_));
 mux2_1 _18429_ (.A0(_03923_),
    .A1(_03926_),
    .S(net793),
    .X(_03927_));
 mux2_1 _18430_ (.A0(net14),
    .A1(_03927_),
    .S(net1498),
    .X(_03928_));
 mux2_1 _18431_ (.A0(\vmem_after_buf[308] ),
    .A1(\vmem_after_buf[292] ),
    .S(net946),
    .X(_03929_));
 mux2_1 _18432_ (.A0(\vmem_after_buf[276] ),
    .A1(\vmem_after_buf[260] ),
    .S(net946),
    .X(_03930_));
 mux2_1 _18433_ (.A0(_03929_),
    .A1(_03930_),
    .S(net909),
    .X(_03931_));
 mux2_1 _18434_ (.A0(\vmem_after_buf[340] ),
    .A1(\vmem_after_buf[324] ),
    .S(net945),
    .X(_03932_));
 mux2_1 _18435_ (.A0(\vmem_after_buf[372] ),
    .A1(\vmem_after_buf[356] ),
    .S(net945),
    .X(_03933_));
 mux2_1 _18436_ (.A0(_03932_),
    .A1(_03933_),
    .S(net904),
    .X(_03934_));
 mux2_1 _18437_ (.A0(_03931_),
    .A1(_03934_),
    .S(net751),
    .X(_03935_));
 mux2_2 _18438_ (.A0(net31),
    .A1(_03935_),
    .S(net1500),
    .X(_03936_));
 a22o_1 _18439_ (.A1(net1478),
    .A2(_03928_),
    .B1(_03936_),
    .B2(net1467),
    .X(_03937_));
 a211o_1 _18440_ (.A1(net1469),
    .A2(_03920_),
    .B1(_03937_),
    .C1(net1471),
    .X(_03938_));
 mux2_1 _18441_ (.A0(\vmem_after_buf[468] ),
    .A1(\vmem_after_buf[452] ),
    .S(net944),
    .X(_03939_));
 mux2_1 _18442_ (.A0(\vmem_after_buf[500] ),
    .A1(\vmem_after_buf[484] ),
    .S(net944),
    .X(_03940_));
 mux2_1 _18443_ (.A0(_03939_),
    .A1(_03940_),
    .S(net902),
    .X(_03941_));
 mux2_1 _18444_ (.A0(\vmem_after_buf[404] ),
    .A1(\vmem_after_buf[388] ),
    .S(net945),
    .X(_03942_));
 mux2_1 _18445_ (.A0(\vmem_after_buf[436] ),
    .A1(\vmem_after_buf[420] ),
    .S(net946),
    .X(_03943_));
 mux2_1 _18446_ (.A0(_03942_),
    .A1(_03943_),
    .S(net902),
    .X(_03944_));
 mux2_1 _18447_ (.A0(_03941_),
    .A1(_03944_),
    .S(net792),
    .X(_03945_));
 mux2_1 _18448_ (.A0(net49),
    .A1(_03945_),
    .S(net1498),
    .X(_03946_));
 o211a_1 _18449_ (.A1(net1470),
    .A2(_03946_),
    .B1(_03938_),
    .C1(net1462),
    .X(_03947_));
 a21o_1 _18450_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[3] ),
    .A2(net1458),
    .B1(net1394),
    .X(_03948_));
 o22a_1 _18451_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[4] ),
    .A2(net1460),
    .B1(_03947_),
    .B2(_03948_),
    .X(_00512_));
 mux2_1 _18452_ (.A0(\vmem_after_buf[341] ),
    .A1(\vmem_after_buf[325] ),
    .S(net920),
    .X(_03949_));
 mux2_1 _18453_ (.A0(\vmem_after_buf[373] ),
    .A1(\vmem_after_buf[357] ),
    .S(net917),
    .X(_03950_));
 mux2_1 _18454_ (.A0(_03949_),
    .A1(_03950_),
    .S(net887),
    .X(_03951_));
 mux2_1 _18455_ (.A0(\vmem_after_buf[277] ),
    .A1(\vmem_after_buf[261] ),
    .S(net917),
    .X(_03952_));
 mux2_1 _18456_ (.A0(\vmem_after_buf[309] ),
    .A1(\vmem_after_buf[293] ),
    .S(net919),
    .X(_03953_));
 mux2_1 _18457_ (.A0(_03952_),
    .A1(_03953_),
    .S(net888),
    .X(_03954_));
 mux2_1 _18458_ (.A0(_03951_),
    .A1(_03954_),
    .S(net760),
    .X(_03955_));
 mux2_1 _18459_ (.A0(net32),
    .A1(_03955_),
    .S(net1494),
    .X(_03956_));
 mux2_1 _18460_ (.A0(\vmem_after_buf[85] ),
    .A1(\vmem_after_buf[69] ),
    .S(net918),
    .X(_03957_));
 mux2_1 _18461_ (.A0(\vmem_after_buf[117] ),
    .A1(\vmem_after_buf[101] ),
    .S(net916),
    .X(_03958_));
 mux2_1 _18462_ (.A0(_03957_),
    .A1(_03958_),
    .S(net887),
    .X(_03959_));
 mux2_1 _18463_ (.A0(\vmem_after_buf[21] ),
    .A1(\vmem_after_buf[5] ),
    .S(net917),
    .X(_03960_));
 mux2_1 _18464_ (.A0(\vmem_after_buf[53] ),
    .A1(\vmem_after_buf[37] ),
    .S(net918),
    .X(_03961_));
 mux2_1 _18465_ (.A0(_03960_),
    .A1(_03961_),
    .S(net887),
    .X(_03962_));
 mux2_1 _18466_ (.A0(_03959_),
    .A1(_03962_),
    .S(net759),
    .X(_03963_));
 mux2_1 _18467_ (.A0(net57),
    .A1(_03963_),
    .S(net1494),
    .X(_03964_));
 mux2_1 _18468_ (.A0(\vmem_after_buf[213] ),
    .A1(\vmem_after_buf[197] ),
    .S(net922),
    .X(_03965_));
 mux2_1 _18469_ (.A0(\vmem_after_buf[245] ),
    .A1(\vmem_after_buf[229] ),
    .S(net918),
    .X(_03966_));
 mux2_1 _18470_ (.A0(_03965_),
    .A1(_03966_),
    .S(net890),
    .X(_03967_));
 mux2_1 _18471_ (.A0(\vmem_after_buf[149] ),
    .A1(\vmem_after_buf[133] ),
    .S(net918),
    .X(_03968_));
 mux2_1 _18472_ (.A0(\vmem_after_buf[181] ),
    .A1(\vmem_after_buf[165] ),
    .S(net918),
    .X(_03969_));
 mux2_1 _18473_ (.A0(_03968_),
    .A1(_03969_),
    .S(net887),
    .X(_03970_));
 mux2_1 _18474_ (.A0(_03967_),
    .A1(_03970_),
    .S(net764),
    .X(_03971_));
 mux2_1 _18475_ (.A0(net15),
    .A1(_03971_),
    .S(net1494),
    .X(_03972_));
 a22o_1 _18476_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[4] ),
    .A2(_03956_),
    .B1(_03972_),
    .B2(net1478),
    .X(_03973_));
 a211o_1 _18477_ (.A1(net1468),
    .A2(_03964_),
    .B1(_03973_),
    .C1(net1472),
    .X(_03974_));
 mux2_1 _18478_ (.A0(\vmem_after_buf[437] ),
    .A1(\vmem_after_buf[421] ),
    .S(net919),
    .X(_03975_));
 mux2_1 _18479_ (.A0(\vmem_after_buf[405] ),
    .A1(\vmem_after_buf[389] ),
    .S(net919),
    .X(_03976_));
 mux2_1 _18480_ (.A0(_03975_),
    .A1(_03976_),
    .S(net906),
    .X(_03977_));
 mux2_1 _18481_ (.A0(\vmem_after_buf[469] ),
    .A1(\vmem_after_buf[453] ),
    .S(net919),
    .X(_03978_));
 mux2_1 _18482_ (.A0(\vmem_after_buf[501] ),
    .A1(\vmem_after_buf[485] ),
    .S(net919),
    .X(_03979_));
 mux2_1 _18483_ (.A0(_03978_),
    .A1(_03979_),
    .S(net889),
    .X(_03980_));
 mux2_1 _18484_ (.A0(_03977_),
    .A1(_03980_),
    .S(net723),
    .X(_03981_));
 mux2_1 _18485_ (.A0(net50),
    .A1(_03981_),
    .S(net1494),
    .X(_03982_));
 or2_1 _18486_ (.A(net1470),
    .B(_03982_),
    .X(_03983_));
 a32o_1 _18487_ (.A1(net1463),
    .A2(_03974_),
    .A3(_03983_),
    .B1(net1458),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[4] ),
    .X(_03984_));
 o22a_1 _18488_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[5] ),
    .A2(net1460),
    .B1(net1394),
    .B2(_03984_),
    .X(_00513_));
 mux2_1 _18489_ (.A0(\vmem_after_buf[54] ),
    .A1(\vmem_after_buf[38] ),
    .S(net949),
    .X(_03985_));
 mux2_1 _18490_ (.A0(\vmem_after_buf[22] ),
    .A1(\vmem_after_buf[6] ),
    .S(net949),
    .X(_03986_));
 mux2_1 _18491_ (.A0(_03985_),
    .A1(_03986_),
    .S(net910),
    .X(_03987_));
 mux2_1 _18492_ (.A0(\vmem_after_buf[86] ),
    .A1(\vmem_after_buf[70] ),
    .S(net949),
    .X(_03988_));
 mux2_1 _18493_ (.A0(\vmem_after_buf[118] ),
    .A1(\vmem_after_buf[102] ),
    .S(net949),
    .X(_03989_));
 mux2_1 _18494_ (.A0(_03988_),
    .A1(_03989_),
    .S(net904),
    .X(_03990_));
 mux2_1 _18495_ (.A0(_03987_),
    .A1(_03990_),
    .S(net754),
    .X(_03991_));
 mux2_2 _18496_ (.A0(net62),
    .A1(_03991_),
    .S(net1499),
    .X(_03992_));
 mux2_1 _18497_ (.A0(\vmem_after_buf[310] ),
    .A1(\vmem_after_buf[294] ),
    .S(net948),
    .X(_03993_));
 mux2_1 _18498_ (.A0(\vmem_after_buf[278] ),
    .A1(\vmem_after_buf[262] ),
    .S(net949),
    .X(_03994_));
 mux2_1 _18499_ (.A0(_03993_),
    .A1(_03994_),
    .S(net911),
    .X(_03995_));
 mux2_1 _18500_ (.A0(\vmem_after_buf[342] ),
    .A1(\vmem_after_buf[326] ),
    .S(net948),
    .X(_03996_));
 mux2_1 _18501_ (.A0(\vmem_after_buf[374] ),
    .A1(\vmem_after_buf[358] ),
    .S(net949),
    .X(_03997_));
 mux2_1 _18502_ (.A0(_03996_),
    .A1(_03997_),
    .S(net903),
    .X(_03998_));
 mux2_1 _18503_ (.A0(_03995_),
    .A1(_03998_),
    .S(net754),
    .X(_03999_));
 mux2_2 _18504_ (.A0(net33),
    .A1(_03999_),
    .S(net1499),
    .X(_04000_));
 mux2_1 _18505_ (.A0(\vmem_after_buf[214] ),
    .A1(\vmem_after_buf[198] ),
    .S(net947),
    .X(_04001_));
 mux2_1 _18506_ (.A0(\vmem_after_buf[246] ),
    .A1(\vmem_after_buf[230] ),
    .S(net948),
    .X(_04002_));
 mux2_1 _18507_ (.A0(_04001_),
    .A1(_04002_),
    .S(net904),
    .X(_04003_));
 mux2_1 _18508_ (.A0(\vmem_after_buf[150] ),
    .A1(\vmem_after_buf[134] ),
    .S(net948),
    .X(_04004_));
 mux2_1 _18509_ (.A0(\vmem_after_buf[182] ),
    .A1(\vmem_after_buf[166] ),
    .S(net948),
    .X(_04005_));
 mux2_1 _18510_ (.A0(_04004_),
    .A1(_04005_),
    .S(net904),
    .X(_04006_));
 mux2_1 _18511_ (.A0(_04003_),
    .A1(_04006_),
    .S(net797),
    .X(_04007_));
 mux2_1 _18512_ (.A0(net16),
    .A1(_04007_),
    .S(net1496),
    .X(_04008_));
 a22o_1 _18513_ (.A1(_03826_),
    .A2(_04000_),
    .B1(_04008_),
    .B2(_03828_),
    .X(_04009_));
 a211o_1 _18514_ (.A1(net1469),
    .A2(_03992_),
    .B1(_04009_),
    .C1(net1472),
    .X(_04010_));
 or2_1 _18515_ (.A(\vmem_after_buf[454] ),
    .B(net954),
    .X(_04011_));
 o211a_1 _18516_ (.A1(\vmem_after_buf[470] ),
    .A2(net948),
    .B1(_04011_),
    .C1(net909),
    .X(_04012_));
 mux2_1 _18517_ (.A0(\vmem_after_buf[502] ),
    .A1(\vmem_after_buf[486] ),
    .S(net948),
    .X(_04013_));
 a211o_1 _18518_ (.A1(net903),
    .A2(_04013_),
    .B1(_04012_),
    .C1(net797),
    .X(_04014_));
 mux2_1 _18519_ (.A0(\vmem_after_buf[406] ),
    .A1(\vmem_after_buf[390] ),
    .S(net948),
    .X(_04015_));
 mux2_1 _18520_ (.A0(\vmem_after_buf[438] ),
    .A1(\vmem_after_buf[422] ),
    .S(net948),
    .X(_04016_));
 mux2_1 _18521_ (.A0(_04015_),
    .A1(_04016_),
    .S(net903),
    .X(_04017_));
 o211a_1 _18522_ (.A1(net755),
    .A2(_04017_),
    .B1(_04014_),
    .C1(net1499),
    .X(_04018_));
 a21oi_2 _18523_ (.A1(net68),
    .A2(net51),
    .B1(_04018_),
    .Y(_04019_));
 nand2_1 _18524_ (.A(net1472),
    .B(_04019_),
    .Y(_04020_));
 a32o_1 _18525_ (.A1(net1463),
    .A2(_04010_),
    .A3(_04020_),
    .B1(net1458),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[5] ),
    .X(_04021_));
 o22a_1 _18526_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[6] ),
    .A2(net1461),
    .B1(net1395),
    .B2(_04021_),
    .X(_00514_));
 mux2_1 _18527_ (.A0(\vmem_after_buf[55] ),
    .A1(\vmem_after_buf[39] ),
    .S(net929),
    .X(_04022_));
 mux2_1 _18528_ (.A0(\vmem_after_buf[23] ),
    .A1(\vmem_after_buf[7] ),
    .S(net927),
    .X(_04023_));
 mux2_1 _18529_ (.A0(_04022_),
    .A1(_04023_),
    .S(net908),
    .X(_04024_));
 mux2_1 _18530_ (.A0(\vmem_after_buf[87] ),
    .A1(\vmem_after_buf[71] ),
    .S(net927),
    .X(_04025_));
 mux2_1 _18531_ (.A0(\vmem_after_buf[119] ),
    .A1(\vmem_after_buf[103] ),
    .S(net929),
    .X(_04026_));
 mux2_1 _18532_ (.A0(_04025_),
    .A1(_04026_),
    .S(net893),
    .X(_04027_));
 mux2_1 _18533_ (.A0(_04024_),
    .A1(_04027_),
    .S(net730),
    .X(_04028_));
 mux2_1 _18534_ (.A0(net63),
    .A1(_04028_),
    .S(net1495),
    .X(_04029_));
 mux2_1 _18535_ (.A0(\vmem_after_buf[183] ),
    .A1(\vmem_after_buf[167] ),
    .S(net929),
    .X(_04030_));
 mux2_1 _18536_ (.A0(\vmem_after_buf[151] ),
    .A1(\vmem_after_buf[135] ),
    .S(net929),
    .X(_04031_));
 mux2_1 _18537_ (.A0(_04030_),
    .A1(_04031_),
    .S(net908),
    .X(_04032_));
 mux2_1 _18538_ (.A0(\vmem_after_buf[215] ),
    .A1(\vmem_after_buf[199] ),
    .S(net930),
    .X(_04033_));
 mux2_1 _18539_ (.A0(\vmem_after_buf[247] ),
    .A1(\vmem_after_buf[231] ),
    .S(net930),
    .X(_04034_));
 mux2_1 _18540_ (.A0(_04033_),
    .A1(_04034_),
    .S(net895),
    .X(_04035_));
 mux2_1 _18541_ (.A0(_04032_),
    .A1(_04035_),
    .S(net733),
    .X(_04036_));
 mux2_1 _18542_ (.A0(net17),
    .A1(_04036_),
    .S(net1495),
    .X(_04037_));
 mux2_1 _18543_ (.A0(\vmem_after_buf[343] ),
    .A1(\vmem_after_buf[327] ),
    .S(net926),
    .X(_04038_));
 mux2_1 _18544_ (.A0(\vmem_after_buf[375] ),
    .A1(\vmem_after_buf[359] ),
    .S(net928),
    .X(_04039_));
 mux2_1 _18545_ (.A0(_04038_),
    .A1(_04039_),
    .S(net893),
    .X(_04040_));
 mux2_1 _18546_ (.A0(\vmem_after_buf[279] ),
    .A1(\vmem_after_buf[263] ),
    .S(net928),
    .X(_04041_));
 mux2_1 _18547_ (.A0(\vmem_after_buf[311] ),
    .A1(\vmem_after_buf[295] ),
    .S(net929),
    .X(_04042_));
 mux2_1 _18548_ (.A0(_04041_),
    .A1(_04042_),
    .S(net893),
    .X(_04043_));
 mux2_1 _18549_ (.A0(_04040_),
    .A1(_04043_),
    .S(net772),
    .X(_04044_));
 mux2_1 _18550_ (.A0(net34),
    .A1(_04044_),
    .S(net1495),
    .X(_04045_));
 a22o_1 _18551_ (.A1(net1468),
    .A2(_04029_),
    .B1(_04045_),
    .B2(net1467),
    .X(_04046_));
 a211o_1 _18552_ (.A1(net1479),
    .A2(_04037_),
    .B1(_04046_),
    .C1(net1471),
    .X(_04047_));
 mux2_1 _18553_ (.A0(\vmem_after_buf[471] ),
    .A1(\vmem_after_buf[455] ),
    .S(net926),
    .X(_04048_));
 mux2_1 _18554_ (.A0(\vmem_after_buf[503] ),
    .A1(\vmem_after_buf[487] ),
    .S(net928),
    .X(_04049_));
 mux2_1 _18555_ (.A0(_04048_),
    .A1(_04049_),
    .S(net893),
    .X(_04050_));
 mux2_1 _18556_ (.A0(\vmem_after_buf[407] ),
    .A1(\vmem_after_buf[391] ),
    .S(net926),
    .X(_04051_));
 mux2_1 _18557_ (.A0(\vmem_after_buf[439] ),
    .A1(\vmem_after_buf[423] ),
    .S(net928),
    .X(_04052_));
 mux2_1 _18558_ (.A0(_04051_),
    .A1(_04052_),
    .S(net894),
    .X(_04053_));
 mux2_1 _18559_ (.A0(_04050_),
    .A1(_04053_),
    .S(net774),
    .X(_04054_));
 mux2_1 _18560_ (.A0(net52),
    .A1(_04054_),
    .S(net1496),
    .X(_04055_));
 or2_1 _18561_ (.A(net1470),
    .B(_04055_),
    .X(_04056_));
 a32o_1 _18562_ (.A1(net1462),
    .A2(_04047_),
    .A3(_04056_),
    .B1(net1459),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[6] ),
    .X(_04057_));
 o22a_1 _18563_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[7] ),
    .A2(net1460),
    .B1(net1394),
    .B2(_04057_),
    .X(_00515_));
 mux2_1 _18564_ (.A0(\vmem_after_buf[88] ),
    .A1(\vmem_after_buf[72] ),
    .S(net921),
    .X(_04058_));
 mux2_1 _18565_ (.A0(\vmem_after_buf[120] ),
    .A1(\vmem_after_buf[104] ),
    .S(net921),
    .X(_04059_));
 mux2_1 _18566_ (.A0(_04058_),
    .A1(_04059_),
    .S(net890),
    .X(_04060_));
 mux2_1 _18567_ (.A0(\vmem_after_buf[24] ),
    .A1(\vmem_after_buf[8] ),
    .S(net921),
    .X(_04061_));
 mux2_1 _18568_ (.A0(\vmem_after_buf[56] ),
    .A1(\vmem_after_buf[40] ),
    .S(net921),
    .X(_04062_));
 mux2_1 _18569_ (.A0(_04061_),
    .A1(_04062_),
    .S(net890),
    .X(_04063_));
 mux2_1 _18570_ (.A0(_04060_),
    .A1(_04063_),
    .S(net765),
    .X(_04064_));
 mux2_1 _18571_ (.A0(net64),
    .A1(_04064_),
    .S(net1492),
    .X(_04065_));
 mux2_1 _18572_ (.A0(\vmem_after_buf[312] ),
    .A1(\vmem_after_buf[296] ),
    .S(net922),
    .X(_04066_));
 mux2_1 _18573_ (.A0(\vmem_after_buf[280] ),
    .A1(\vmem_after_buf[264] ),
    .S(net922),
    .X(_04067_));
 mux2_1 _18574_ (.A0(_04066_),
    .A1(_04067_),
    .S(net906),
    .X(_04068_));
 mux2_1 _18575_ (.A0(\vmem_after_buf[344] ),
    .A1(\vmem_after_buf[328] ),
    .S(net921),
    .X(_04069_));
 mux2_1 _18576_ (.A0(\vmem_after_buf[376] ),
    .A1(\vmem_after_buf[360] ),
    .S(net922),
    .X(_04070_));
 mux2_1 _18577_ (.A0(_04069_),
    .A1(_04070_),
    .S(net890),
    .X(_04071_));
 mux2_1 _18578_ (.A0(_04068_),
    .A1(_04071_),
    .S(net725),
    .X(_04072_));
 mux2_1 _18579_ (.A0(net36),
    .A1(_04072_),
    .S(net1492),
    .X(_04073_));
 mux2_1 _18580_ (.A0(\vmem_after_buf[216] ),
    .A1(\vmem_after_buf[200] ),
    .S(net920),
    .X(_04074_));
 mux2_1 _18581_ (.A0(\vmem_after_buf[248] ),
    .A1(\vmem_after_buf[232] ),
    .S(net920),
    .X(_04075_));
 mux2_1 _18582_ (.A0(_04074_),
    .A1(_04075_),
    .S(net890),
    .X(_04076_));
 mux2_1 _18583_ (.A0(\vmem_after_buf[152] ),
    .A1(\vmem_after_buf[136] ),
    .S(net920),
    .X(_04077_));
 mux2_1 _18584_ (.A0(\vmem_after_buf[184] ),
    .A1(\vmem_after_buf[168] ),
    .S(net920),
    .X(_04078_));
 mux2_1 _18585_ (.A0(_04077_),
    .A1(_04078_),
    .S(net890),
    .X(_04079_));
 mux2_1 _18586_ (.A0(_04076_),
    .A1(_04079_),
    .S(net763),
    .X(_04080_));
 mux2_1 _18587_ (.A0(net18),
    .A1(_04080_),
    .S(net1492),
    .X(_04081_));
 a22o_1 _18588_ (.A1(net1467),
    .A2(_04073_),
    .B1(_04081_),
    .B2(_03828_),
    .X(_04082_));
 a211o_1 _18589_ (.A1(net1468),
    .A2(_04065_),
    .B1(_04082_),
    .C1(net1472),
    .X(_04083_));
 mux2_1 _18590_ (.A0(\vmem_after_buf[472] ),
    .A1(\vmem_after_buf[456] ),
    .S(net920),
    .X(_04084_));
 mux2_1 _18591_ (.A0(\vmem_after_buf[504] ),
    .A1(\vmem_after_buf[488] ),
    .S(net920),
    .X(_04085_));
 mux2_1 _18592_ (.A0(_04084_),
    .A1(_04085_),
    .S(net890),
    .X(_04086_));
 mux2_1 _18593_ (.A0(\vmem_after_buf[408] ),
    .A1(\vmem_after_buf[392] ),
    .S(net920),
    .X(_04087_));
 mux2_1 _18594_ (.A0(\vmem_after_buf[440] ),
    .A1(\vmem_after_buf[424] ),
    .S(net920),
    .X(_04088_));
 mux2_1 _18595_ (.A0(_04087_),
    .A1(_04088_),
    .S(net890),
    .X(_04089_));
 mux2_1 _18596_ (.A0(_04086_),
    .A1(_04089_),
    .S(net764),
    .X(_04090_));
 mux2_1 _18597_ (.A0(net53),
    .A1(_04090_),
    .S(net1492),
    .X(_04091_));
 o211a_1 _18598_ (.A1(net1470),
    .A2(_04091_),
    .B1(_04083_),
    .C1(net1462),
    .X(_04092_));
 a21o_1 _18599_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[7] ),
    .A2(net1458),
    .B1(net1394),
    .X(_04093_));
 o22a_1 _18600_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[8] ),
    .A2(net1460),
    .B1(_04092_),
    .B2(_04093_),
    .X(_00516_));
 mux2_1 _18601_ (.A0(\vmem_after_buf[89] ),
    .A1(\vmem_after_buf[73] ),
    .S(net924),
    .X(_04094_));
 mux2_1 _18602_ (.A0(\vmem_after_buf[121] ),
    .A1(\vmem_after_buf[105] ),
    .S(net924),
    .X(_04095_));
 mux2_1 _18603_ (.A0(_04094_),
    .A1(_04095_),
    .S(_03760_),
    .X(_04096_));
 mux2_1 _18604_ (.A0(\vmem_after_buf[25] ),
    .A1(\vmem_after_buf[9] ),
    .S(net924),
    .X(_04097_));
 mux2_1 _18605_ (.A0(\vmem_after_buf[57] ),
    .A1(\vmem_after_buf[41] ),
    .S(net939),
    .X(_04098_));
 mux2_1 _18606_ (.A0(_04097_),
    .A1(_04098_),
    .S(_03760_),
    .X(_04099_));
 mux2_1 _18607_ (.A0(_04096_),
    .A1(_04099_),
    .S(net769),
    .X(_04100_));
 mux2_1 _18608_ (.A0(net65),
    .A1(_04100_),
    .S(net1493),
    .X(_04101_));
 mux2_1 _18609_ (.A0(\vmem_after_buf[345] ),
    .A1(\vmem_after_buf[329] ),
    .S(net929),
    .X(_04102_));
 mux2_1 _18610_ (.A0(\vmem_after_buf[377] ),
    .A1(\vmem_after_buf[361] ),
    .S(net939),
    .X(_04103_));
 mux2_1 _18611_ (.A0(_04102_),
    .A1(_04103_),
    .S(net895),
    .X(_04104_));
 mux2_1 _18612_ (.A0(\vmem_after_buf[281] ),
    .A1(\vmem_after_buf[265] ),
    .S(net929),
    .X(_04105_));
 mux2_1 _18613_ (.A0(\vmem_after_buf[313] ),
    .A1(\vmem_after_buf[297] ),
    .S(net939),
    .X(_04106_));
 mux2_1 _18614_ (.A0(_04105_),
    .A1(_04106_),
    .S(net900),
    .X(_04107_));
 mux2_1 _18615_ (.A0(_04104_),
    .A1(_04107_),
    .S(net786),
    .X(_04108_));
 mux2_1 _18616_ (.A0(net37),
    .A1(_04108_),
    .S(net1493),
    .X(_04109_));
 mux2_1 _18617_ (.A0(\vmem_after_buf[217] ),
    .A1(\vmem_after_buf[201] ),
    .S(net929),
    .X(_04110_));
 mux2_1 _18618_ (.A0(\vmem_after_buf[249] ),
    .A1(\vmem_after_buf[233] ),
    .S(net939),
    .X(_04111_));
 mux2_1 _18619_ (.A0(_04110_),
    .A1(_04111_),
    .S(net891),
    .X(_04112_));
 mux2_1 _18620_ (.A0(\vmem_after_buf[153] ),
    .A1(\vmem_after_buf[137] ),
    .S(net923),
    .X(_04113_));
 mux2_1 _18621_ (.A0(\vmem_after_buf[185] ),
    .A1(\vmem_after_buf[169] ),
    .S(net939),
    .X(_04114_));
 mux2_1 _18622_ (.A0(_04113_),
    .A1(_04114_),
    .S(net892),
    .X(_04115_));
 mux2_1 _18623_ (.A0(_04112_),
    .A1(_04115_),
    .S(net767),
    .X(_04116_));
 mux2_1 _18624_ (.A0(net19),
    .A1(_04116_),
    .S(net1492),
    .X(_04117_));
 a22o_1 _18625_ (.A1(_03826_),
    .A2(_04109_),
    .B1(_04117_),
    .B2(_03828_),
    .X(_04118_));
 a211o_1 _18626_ (.A1(net1468),
    .A2(_04101_),
    .B1(_04118_),
    .C1(net1472),
    .X(_04119_));
 mux2_1 _18627_ (.A0(\vmem_after_buf[473] ),
    .A1(\vmem_after_buf[457] ),
    .S(net939),
    .X(_04120_));
 mux2_1 _18628_ (.A0(\vmem_after_buf[505] ),
    .A1(\vmem_after_buf[489] ),
    .S(net941),
    .X(_04121_));
 mux2_1 _18629_ (.A0(_04120_),
    .A1(_04121_),
    .S(net900),
    .X(_04122_));
 mux2_1 _18630_ (.A0(\vmem_after_buf[409] ),
    .A1(\vmem_after_buf[393] ),
    .S(net939),
    .X(_04123_));
 mux2_1 _18631_ (.A0(\vmem_after_buf[441] ),
    .A1(\vmem_after_buf[425] ),
    .S(net939),
    .X(_04124_));
 mux2_1 _18632_ (.A0(_04123_),
    .A1(_04124_),
    .S(net900),
    .X(_04125_));
 mux2_1 _18633_ (.A0(_04122_),
    .A1(_04125_),
    .S(net788),
    .X(_04126_));
 mux2_1 _18634_ (.A0(net54),
    .A1(_04126_),
    .S(net1499),
    .X(_04127_));
 o211a_1 _18635_ (.A1(_03758_),
    .A2(_04127_),
    .B1(_04119_),
    .C1(net1463),
    .X(_04128_));
 a21o_1 _18636_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[8] ),
    .A2(net1458),
    .B1(net1394),
    .X(_04129_));
 o22a_1 _18637_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[9] ),
    .A2(net1460),
    .B1(_04128_),
    .B2(_04129_),
    .X(_00517_));
 mux2_1 _18638_ (.A0(\vmem_after_buf[90] ),
    .A1(\vmem_after_buf[74] ),
    .S(net927),
    .X(_04130_));
 mux2_1 _18639_ (.A0(\vmem_after_buf[122] ),
    .A1(\vmem_after_buf[106] ),
    .S(net927),
    .X(_04131_));
 mux2_1 _18640_ (.A0(_04130_),
    .A1(_04131_),
    .S(net893),
    .X(_04132_));
 mux2_1 _18641_ (.A0(\vmem_after_buf[26] ),
    .A1(\vmem_after_buf[10] ),
    .S(net927),
    .X(_04133_));
 mux2_1 _18642_ (.A0(\vmem_after_buf[58] ),
    .A1(\vmem_after_buf[42] ),
    .S(net927),
    .X(_04134_));
 mux2_1 _18643_ (.A0(_04133_),
    .A1(_04134_),
    .S(net893),
    .X(_04135_));
 mux2_1 _18644_ (.A0(_04132_),
    .A1(_04135_),
    .S(net770),
    .X(_04136_));
 mux2_1 _18645_ (.A0(net3),
    .A1(_04136_),
    .S(net1495),
    .X(_04137_));
 mux2_1 _18646_ (.A0(\vmem_after_buf[346] ),
    .A1(\vmem_after_buf[330] ),
    .S(net925),
    .X(_04138_));
 mux2_1 _18647_ (.A0(\vmem_after_buf[378] ),
    .A1(\vmem_after_buf[362] ),
    .S(net925),
    .X(_04139_));
 mux2_1 _18648_ (.A0(_04138_),
    .A1(_04139_),
    .S(net894),
    .X(_04140_));
 mux2_1 _18649_ (.A0(\vmem_after_buf[282] ),
    .A1(\vmem_after_buf[266] ),
    .S(net925),
    .X(_04141_));
 mux2_1 _18650_ (.A0(\vmem_after_buf[314] ),
    .A1(\vmem_after_buf[298] ),
    .S(net925),
    .X(_04142_));
 mux2_1 _18651_ (.A0(_04141_),
    .A1(_04142_),
    .S(net894),
    .X(_04143_));
 mux2_1 _18652_ (.A0(_04140_),
    .A1(_04143_),
    .S(net772),
    .X(_04144_));
 mux2_1 _18653_ (.A0(net38),
    .A1(_04144_),
    .S(net1495),
    .X(_04145_));
 mux2_1 _18654_ (.A0(\vmem_after_buf[186] ),
    .A1(\vmem_after_buf[170] ),
    .S(net921),
    .X(_04146_));
 mux2_1 _18655_ (.A0(\vmem_after_buf[154] ),
    .A1(\vmem_after_buf[138] ),
    .S(net927),
    .X(_04147_));
 mux2_1 _18656_ (.A0(_04146_),
    .A1(_04147_),
    .S(_03759_),
    .X(_04148_));
 mux2_1 _18657_ (.A0(\vmem_after_buf[218] ),
    .A1(\vmem_after_buf[202] ),
    .S(net921),
    .X(_04149_));
 mux2_1 _18658_ (.A0(\vmem_after_buf[250] ),
    .A1(\vmem_after_buf[234] ),
    .S(net921),
    .X(_04150_));
 mux2_1 _18659_ (.A0(_04149_),
    .A1(_04150_),
    .S(net891),
    .X(_04151_));
 mux2_1 _18660_ (.A0(_04148_),
    .A1(_04151_),
    .S(net725),
    .X(_04152_));
 mux2_1 _18661_ (.A0(net20),
    .A1(_04152_),
    .S(net1492),
    .X(_04153_));
 a22o_1 _18662_ (.A1(net1467),
    .A2(_04145_),
    .B1(_04153_),
    .B2(_03828_),
    .X(_04154_));
 a211o_1 _18663_ (.A1(net1468),
    .A2(_04137_),
    .B1(_04154_),
    .C1(net1472),
    .X(_04155_));
 mux2_1 _18664_ (.A0(\vmem_after_buf[474] ),
    .A1(\vmem_after_buf[458] ),
    .S(net927),
    .X(_04156_));
 mux2_1 _18665_ (.A0(\vmem_after_buf[506] ),
    .A1(\vmem_after_buf[490] ),
    .S(net927),
    .X(_04157_));
 mux2_1 _18666_ (.A0(_04156_),
    .A1(_04157_),
    .S(net893),
    .X(_04158_));
 mux2_1 _18667_ (.A0(\vmem_after_buf[410] ),
    .A1(\vmem_after_buf[394] ),
    .S(net921),
    .X(_04159_));
 mux2_1 _18668_ (.A0(\vmem_after_buf[442] ),
    .A1(\vmem_after_buf[426] ),
    .S(net921),
    .X(_04160_));
 mux2_1 _18669_ (.A0(_04159_),
    .A1(_04160_),
    .S(net891),
    .X(_04161_));
 mux2_1 _18670_ (.A0(_04158_),
    .A1(_04161_),
    .S(net765),
    .X(_04162_));
 mux2_1 _18671_ (.A0(net55),
    .A1(_04162_),
    .S(net1492),
    .X(_04163_));
 o211a_1 _18672_ (.A1(net1470),
    .A2(_04163_),
    .B1(_04155_),
    .C1(net1462),
    .X(_04164_));
 a21o_1 _18673_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[9] ),
    .A2(net1458),
    .B1(net1394),
    .X(_04165_));
 o22a_1 _18674_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[10] ),
    .A2(net1460),
    .B1(_04164_),
    .B2(_04165_),
    .X(_00518_));
 mux2_1 _18675_ (.A0(\vmem_after_buf[91] ),
    .A1(\vmem_after_buf[75] ),
    .S(net932),
    .X(_04166_));
 mux2_1 _18676_ (.A0(\vmem_after_buf[123] ),
    .A1(\vmem_after_buf[107] ),
    .S(net932),
    .X(_04167_));
 mux2_1 _18677_ (.A0(_04166_),
    .A1(_04167_),
    .S(net899),
    .X(_04168_));
 mux2_1 _18678_ (.A0(\vmem_after_buf[27] ),
    .A1(\vmem_after_buf[11] ),
    .S(net932),
    .X(_04169_));
 mux2_1 _18679_ (.A0(\vmem_after_buf[59] ),
    .A1(\vmem_after_buf[43] ),
    .S(net932),
    .X(_04170_));
 mux2_1 _18680_ (.A0(_04169_),
    .A1(_04170_),
    .S(net899),
    .X(_04171_));
 mux2_1 _18681_ (.A0(_04168_),
    .A1(_04171_),
    .S(net779),
    .X(_04172_));
 mux2_2 _18682_ (.A0(net4),
    .A1(_04172_),
    .S(net1497),
    .X(_04173_));
 mux2_1 _18683_ (.A0(\vmem_after_buf[187] ),
    .A1(\vmem_after_buf[171] ),
    .S(net933),
    .X(_04174_));
 mux2_1 _18684_ (.A0(\vmem_after_buf[155] ),
    .A1(\vmem_after_buf[139] ),
    .S(net931),
    .X(_04175_));
 mux2_1 _18685_ (.A0(_04174_),
    .A1(_04175_),
    .S(net907),
    .X(_04176_));
 mux2_1 _18686_ (.A0(\vmem_after_buf[219] ),
    .A1(\vmem_after_buf[203] ),
    .S(net938),
    .X(_04177_));
 mux2_1 _18687_ (.A0(\vmem_after_buf[251] ),
    .A1(\vmem_after_buf[235] ),
    .S(net933),
    .X(_04178_));
 mux2_1 _18688_ (.A0(_04177_),
    .A1(_04178_),
    .S(net896),
    .X(_04179_));
 mux2_1 _18689_ (.A0(_04176_),
    .A1(_04179_),
    .S(net738),
    .X(_04180_));
 mux2_1 _18690_ (.A0(net21),
    .A1(_04180_),
    .S(net1495),
    .X(_04181_));
 mux2_1 _18691_ (.A0(\vmem_after_buf[315] ),
    .A1(\vmem_after_buf[299] ),
    .S(net932),
    .X(_04182_));
 mux2_1 _18692_ (.A0(\vmem_after_buf[283] ),
    .A1(\vmem_after_buf[267] ),
    .S(net932),
    .X(_04183_));
 mux2_1 _18693_ (.A0(_04182_),
    .A1(_04183_),
    .S(net907),
    .X(_04184_));
 mux2_1 _18694_ (.A0(\vmem_after_buf[347] ),
    .A1(\vmem_after_buf[331] ),
    .S(net932),
    .X(_04185_));
 mux2_1 _18695_ (.A0(\vmem_after_buf[379] ),
    .A1(\vmem_after_buf[363] ),
    .S(net932),
    .X(_04186_));
 mux2_1 _18696_ (.A0(_04185_),
    .A1(_04186_),
    .S(net896),
    .X(_04187_));
 mux2_1 _18697_ (.A0(_04184_),
    .A1(_04187_),
    .S(net737),
    .X(_04188_));
 mux2_2 _18698_ (.A0(net39),
    .A1(_04188_),
    .S(net1497),
    .X(_04189_));
 a22o_1 _18699_ (.A1(net1468),
    .A2(_04173_),
    .B1(_04181_),
    .B2(net1479),
    .X(_04190_));
 a211o_1 _18700_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[4] ),
    .A2(_04189_),
    .B1(_04190_),
    .C1(net1471),
    .X(_04191_));
 mux2_1 _18701_ (.A0(\vmem_after_buf[475] ),
    .A1(\vmem_after_buf[459] ),
    .S(net932),
    .X(_04192_));
 mux2_1 _18702_ (.A0(\vmem_after_buf[507] ),
    .A1(\vmem_after_buf[491] ),
    .S(net933),
    .X(_04193_));
 mux2_1 _18703_ (.A0(_04192_),
    .A1(_04193_),
    .S(net896),
    .X(_04194_));
 mux2_1 _18704_ (.A0(\vmem_after_buf[411] ),
    .A1(\vmem_after_buf[395] ),
    .S(net933),
    .X(_04195_));
 mux2_1 _18705_ (.A0(\vmem_after_buf[443] ),
    .A1(\vmem_after_buf[427] ),
    .S(net933),
    .X(_04196_));
 mux2_1 _18706_ (.A0(_04195_),
    .A1(_04196_),
    .S(net899),
    .X(_04197_));
 mux2_1 _18707_ (.A0(_04194_),
    .A1(_04197_),
    .S(net780),
    .X(_04198_));
 mux2_1 _18708_ (.A0(net56),
    .A1(_04198_),
    .S(net1497),
    .X(_04199_));
 o211a_1 _18709_ (.A1(net1470),
    .A2(_04199_),
    .B1(_04191_),
    .C1(net1462),
    .X(_04200_));
 a21o_1 _18710_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[10] ),
    .A2(net1458),
    .B1(net1394),
    .X(_04201_));
 o22a_1 _18711_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[11] ),
    .A2(net1460),
    .B1(_04200_),
    .B2(_04201_),
    .X(_00519_));
 mux2_1 _18712_ (.A0(\vmem_after_buf[92] ),
    .A1(\vmem_after_buf[76] ),
    .S(net947),
    .X(_04202_));
 mux2_1 _18713_ (.A0(\vmem_after_buf[124] ),
    .A1(\vmem_after_buf[108] ),
    .S(net943),
    .X(_04203_));
 mux2_1 _18714_ (.A0(_04202_),
    .A1(_04203_),
    .S(net901),
    .X(_04204_));
 mux2_1 _18715_ (.A0(\vmem_after_buf[28] ),
    .A1(\vmem_after_buf[12] ),
    .S(net942),
    .X(_04205_));
 mux2_1 _18716_ (.A0(\vmem_after_buf[60] ),
    .A1(\vmem_after_buf[44] ),
    .S(net943),
    .X(_04206_));
 mux2_1 _18717_ (.A0(_04205_),
    .A1(_04206_),
    .S(net905),
    .X(_04207_));
 mux2_1 _18718_ (.A0(_04204_),
    .A1(_04207_),
    .S(net790),
    .X(_04208_));
 mux2_2 _18719_ (.A0(net5),
    .A1(_04208_),
    .S(net1499),
    .X(_04209_));
 mux2_1 _18720_ (.A0(\vmem_after_buf[348] ),
    .A1(\vmem_after_buf[332] ),
    .S(net947),
    .X(_04210_));
 mux2_1 _18721_ (.A0(\vmem_after_buf[380] ),
    .A1(\vmem_after_buf[364] ),
    .S(net947),
    .X(_04211_));
 mux2_1 _18722_ (.A0(_04210_),
    .A1(_04211_),
    .S(net903),
    .X(_04212_));
 mux2_1 _18723_ (.A0(\vmem_after_buf[284] ),
    .A1(\vmem_after_buf[268] ),
    .S(net950),
    .X(_04213_));
 mux2_1 _18724_ (.A0(\vmem_after_buf[316] ),
    .A1(\vmem_after_buf[300] ),
    .S(net950),
    .X(_04214_));
 mux2_1 _18725_ (.A0(_04213_),
    .A1(_04214_),
    .S(net903),
    .X(_04215_));
 mux2_1 _18726_ (.A0(_04212_),
    .A1(_04215_),
    .S(net799),
    .X(_04216_));
 mux2_2 _18727_ (.A0(net40),
    .A1(_04216_),
    .S(net1499),
    .X(_04217_));
 mux2_1 _18728_ (.A0(\vmem_after_buf[188] ),
    .A1(\vmem_after_buf[172] ),
    .S(net942),
    .X(_04218_));
 mux2_1 _18729_ (.A0(\vmem_after_buf[156] ),
    .A1(\vmem_after_buf[140] ),
    .S(net947),
    .X(_04219_));
 mux2_1 _18730_ (.A0(_04218_),
    .A1(_04219_),
    .S(net910),
    .X(_04220_));
 mux2_1 _18731_ (.A0(\vmem_after_buf[220] ),
    .A1(\vmem_after_buf[204] ),
    .S(net947),
    .X(_04221_));
 mux2_1 _18732_ (.A0(\vmem_after_buf[252] ),
    .A1(\vmem_after_buf[236] ),
    .S(net942),
    .X(_04222_));
 mux2_1 _18733_ (.A0(_04221_),
    .A1(_04222_),
    .S(net901),
    .X(_04223_));
 mux2_1 _18734_ (.A0(_04220_),
    .A1(_04223_),
    .S(net746),
    .X(_04224_));
 mux2_1 _18735_ (.A0(net22),
    .A1(_04224_),
    .S(net1496),
    .X(_04225_));
 a22o_1 _18736_ (.A1(net1467),
    .A2(_04217_),
    .B1(_04225_),
    .B2(_03828_),
    .X(_04226_));
 a211o_1 _18737_ (.A1(net1469),
    .A2(_04209_),
    .B1(_04226_),
    .C1(net1471),
    .X(_04227_));
 mux2_1 _18738_ (.A0(\vmem_after_buf[444] ),
    .A1(\vmem_after_buf[428] ),
    .S(net947),
    .X(_04228_));
 mux2_1 _18739_ (.A0(\vmem_after_buf[412] ),
    .A1(\vmem_after_buf[396] ),
    .S(net947),
    .X(_04229_));
 mux2_1 _18740_ (.A0(_04228_),
    .A1(_04229_),
    .S(net911),
    .X(_04230_));
 mux2_1 _18741_ (.A0(\vmem_after_buf[476] ),
    .A1(\vmem_after_buf[460] ),
    .S(net947),
    .X(_04231_));
 mux2_1 _18742_ (.A0(\vmem_after_buf[508] ),
    .A1(\vmem_after_buf[492] ),
    .S(net947),
    .X(_04232_));
 mux2_1 _18743_ (.A0(_04231_),
    .A1(_04232_),
    .S(net903),
    .X(_04233_));
 mux2_1 _18744_ (.A0(_04230_),
    .A1(_04233_),
    .S(net753),
    .X(_04234_));
 mux2_2 _18745_ (.A0(net58),
    .A1(_04234_),
    .S(net1499),
    .X(_04235_));
 o211a_1 _18746_ (.A1(net1470),
    .A2(_04235_),
    .B1(_04227_),
    .C1(net1463),
    .X(_04236_));
 a21o_1 _18747_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[11] ),
    .A2(net1458),
    .B1(net1395),
    .X(_04237_));
 o22a_1 _18748_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[12] ),
    .A2(net1461),
    .B1(_04236_),
    .B2(_04237_),
    .X(_00520_));
 mux2_1 _18749_ (.A0(\vmem_after_buf[93] ),
    .A1(\vmem_after_buf[77] ),
    .S(net928),
    .X(_04238_));
 mux2_1 _18750_ (.A0(\vmem_after_buf[125] ),
    .A1(\vmem_after_buf[109] ),
    .S(net928),
    .X(_04239_));
 mux2_1 _18751_ (.A0(_04238_),
    .A1(_04239_),
    .S(net895),
    .X(_04240_));
 mux2_1 _18752_ (.A0(\vmem_after_buf[29] ),
    .A1(\vmem_after_buf[13] ),
    .S(net928),
    .X(_04241_));
 mux2_1 _18753_ (.A0(\vmem_after_buf[61] ),
    .A1(\vmem_after_buf[45] ),
    .S(net934),
    .X(_04242_));
 mux2_1 _18754_ (.A0(_04241_),
    .A1(_04242_),
    .S(net895),
    .X(_04243_));
 mux2_1 _18755_ (.A0(_04240_),
    .A1(_04243_),
    .S(net774),
    .X(_04244_));
 mux2_1 _18756_ (.A0(net6),
    .A1(_04244_),
    .S(net1496),
    .X(_04245_));
 mux2_1 _18757_ (.A0(\vmem_after_buf[349] ),
    .A1(\vmem_after_buf[333] ),
    .S(net934),
    .X(_04246_));
 mux2_1 _18758_ (.A0(\vmem_after_buf[381] ),
    .A1(\vmem_after_buf[365] ),
    .S(net934),
    .X(_04247_));
 mux2_1 _18759_ (.A0(_04246_),
    .A1(_04247_),
    .S(net897),
    .X(_04248_));
 mux2_1 _18760_ (.A0(\vmem_after_buf[285] ),
    .A1(\vmem_after_buf[269] ),
    .S(net934),
    .X(_04249_));
 mux2_1 _18761_ (.A0(\vmem_after_buf[317] ),
    .A1(\vmem_after_buf[301] ),
    .S(net934),
    .X(_04250_));
 mux2_1 _18762_ (.A0(_04249_),
    .A1(_04250_),
    .S(net897),
    .X(_04251_));
 mux2_1 _18763_ (.A0(_04248_),
    .A1(_04251_),
    .S(net781),
    .X(_04252_));
 mux2_1 _18764_ (.A0(net41),
    .A1(_04252_),
    .S(net1497),
    .X(_04253_));
 mux2_1 _18765_ (.A0(\vmem_after_buf[221] ),
    .A1(\vmem_after_buf[205] ),
    .S(net937),
    .X(_04254_));
 mux2_1 _18766_ (.A0(\vmem_after_buf[253] ),
    .A1(\vmem_after_buf[237] ),
    .S(net937),
    .X(_04255_));
 mux2_1 _18767_ (.A0(_04254_),
    .A1(_04255_),
    .S(net897),
    .X(_04256_));
 mux2_1 _18768_ (.A0(\vmem_after_buf[157] ),
    .A1(\vmem_after_buf[141] ),
    .S(net934),
    .X(_04257_));
 mux2_1 _18769_ (.A0(\vmem_after_buf[189] ),
    .A1(\vmem_after_buf[173] ),
    .S(net934),
    .X(_04258_));
 mux2_1 _18770_ (.A0(_04257_),
    .A1(_04258_),
    .S(net897),
    .X(_04259_));
 mux2_1 _18771_ (.A0(_04256_),
    .A1(_04259_),
    .S(net781),
    .X(_04260_));
 mux2_1 _18772_ (.A0(net23),
    .A1(_04260_),
    .S(net1497),
    .X(_04261_));
 a22o_1 _18773_ (.A1(net1467),
    .A2(_04253_),
    .B1(_04261_),
    .B2(_03828_),
    .X(_04262_));
 a211o_1 _18774_ (.A1(net1469),
    .A2(_04245_),
    .B1(_04262_),
    .C1(net1472),
    .X(_04263_));
 mux2_1 _18775_ (.A0(\vmem_after_buf[445] ),
    .A1(\vmem_after_buf[429] ),
    .S(net934),
    .X(_04264_));
 mux2_1 _18776_ (.A0(\vmem_after_buf[413] ),
    .A1(\vmem_after_buf[397] ),
    .S(net928),
    .X(_04265_));
 mux2_1 _18777_ (.A0(_04264_),
    .A1(_04265_),
    .S(net908),
    .X(_04266_));
 mux2_1 _18778_ (.A0(\vmem_after_buf[477] ),
    .A1(\vmem_after_buf[461] ),
    .S(net929),
    .X(_04267_));
 mux2_1 _18779_ (.A0(\vmem_after_buf[509] ),
    .A1(\vmem_after_buf[493] ),
    .S(net928),
    .X(_04268_));
 mux2_1 _18780_ (.A0(_04267_),
    .A1(_04268_),
    .S(net895),
    .X(_04269_));
 mux2_1 _18781_ (.A0(_04266_),
    .A1(_04269_),
    .S(net734),
    .X(_04270_));
 mux2_1 _18782_ (.A0(net59),
    .A1(_04270_),
    .S(net1495),
    .X(_04271_));
 o211a_1 _18783_ (.A1(net1470),
    .A2(_04271_),
    .B1(_04263_),
    .C1(net1462),
    .X(_04272_));
 a21o_1 _18784_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[12] ),
    .A2(net1459),
    .B1(net1395),
    .X(_04273_));
 o22a_1 _18785_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[13] ),
    .A2(net1461),
    .B1(_04272_),
    .B2(_04273_),
    .X(_00521_));
 mux2_1 _18786_ (.A0(\vmem_after_buf[94] ),
    .A1(\vmem_after_buf[78] ),
    .S(net935),
    .X(_04274_));
 mux2_1 _18787_ (.A0(\vmem_after_buf[126] ),
    .A1(\vmem_after_buf[110] ),
    .S(net935),
    .X(_04275_));
 mux2_1 _18788_ (.A0(_04274_),
    .A1(_04275_),
    .S(net897),
    .X(_04276_));
 mux2_1 _18789_ (.A0(\vmem_after_buf[30] ),
    .A1(\vmem_after_buf[14] ),
    .S(net935),
    .X(_04277_));
 mux2_1 _18790_ (.A0(\vmem_after_buf[62] ),
    .A1(\vmem_after_buf[46] ),
    .S(net936),
    .X(_04278_));
 mux2_1 _18791_ (.A0(_04277_),
    .A1(_04278_),
    .S(net897),
    .X(_04279_));
 mux2_1 _18792_ (.A0(_04276_),
    .A1(_04279_),
    .S(net782),
    .X(_04280_));
 mux2_1 _18793_ (.A0(net7),
    .A1(_04280_),
    .S(net1497),
    .X(_04281_));
 mux2_1 _18794_ (.A0(\vmem_after_buf[350] ),
    .A1(\vmem_after_buf[334] ),
    .S(net935),
    .X(_04282_));
 mux2_1 _18795_ (.A0(\vmem_after_buf[382] ),
    .A1(\vmem_after_buf[366] ),
    .S(net935),
    .X(_04283_));
 mux2_1 _18796_ (.A0(_04282_),
    .A1(_04283_),
    .S(net898),
    .X(_04284_));
 mux2_1 _18797_ (.A0(\vmem_after_buf[286] ),
    .A1(\vmem_after_buf[270] ),
    .S(net935),
    .X(_04285_));
 mux2_1 _18798_ (.A0(\vmem_after_buf[318] ),
    .A1(\vmem_after_buf[302] ),
    .S(net935),
    .X(_04286_));
 mux2_1 _18799_ (.A0(_04285_),
    .A1(_04286_),
    .S(net898),
    .X(_04287_));
 mux2_1 _18800_ (.A0(_04284_),
    .A1(_04287_),
    .S(net782),
    .X(_04288_));
 mux2_1 _18801_ (.A0(net42),
    .A1(_04288_),
    .S(net1497),
    .X(_04289_));
 mux2_1 _18802_ (.A0(\vmem_after_buf[222] ),
    .A1(\vmem_after_buf[206] ),
    .S(net934),
    .X(_04290_));
 mux2_1 _18803_ (.A0(\vmem_after_buf[254] ),
    .A1(\vmem_after_buf[238] ),
    .S(net936),
    .X(_04291_));
 mux2_1 _18804_ (.A0(_04290_),
    .A1(_04291_),
    .S(net897),
    .X(_04292_));
 mux2_1 _18805_ (.A0(\vmem_after_buf[158] ),
    .A1(\vmem_after_buf[142] ),
    .S(net936),
    .X(_04293_));
 mux2_1 _18806_ (.A0(\vmem_after_buf[190] ),
    .A1(\vmem_after_buf[174] ),
    .S(net936),
    .X(_04294_));
 mux2_1 _18807_ (.A0(_04293_),
    .A1(_04294_),
    .S(net897),
    .X(_04295_));
 mux2_1 _18808_ (.A0(_04292_),
    .A1(_04295_),
    .S(net781),
    .X(_04296_));
 mux2_1 _18809_ (.A0(net25),
    .A1(_04296_),
    .S(net1496),
    .X(_04297_));
 a22o_1 _18810_ (.A1(net1467),
    .A2(_04289_),
    .B1(_04297_),
    .B2(_03828_),
    .X(_04298_));
 a211o_1 _18811_ (.A1(net1468),
    .A2(_04281_),
    .B1(_04298_),
    .C1(net1471),
    .X(_04299_));
 or2_1 _18812_ (.A(\vmem_after_buf[462] ),
    .B(net953),
    .X(_04300_));
 o211a_1 _18813_ (.A1(\vmem_after_buf[478] ),
    .A2(net935),
    .B1(_04300_),
    .C1(net911),
    .X(_04301_));
 mux2_1 _18814_ (.A0(\vmem_after_buf[510] ),
    .A1(\vmem_after_buf[494] ),
    .S(net935),
    .X(_04302_));
 a211o_1 _18815_ (.A1(net898),
    .A2(_04302_),
    .B1(_04301_),
    .C1(net783),
    .X(_04303_));
 mux2_1 _18816_ (.A0(\vmem_after_buf[414] ),
    .A1(\vmem_after_buf[398] ),
    .S(net936),
    .X(_04304_));
 mux2_1 _18817_ (.A0(\vmem_after_buf[446] ),
    .A1(\vmem_after_buf[430] ),
    .S(net936),
    .X(_04305_));
 mux2_1 _18818_ (.A0(_04304_),
    .A1(_04305_),
    .S(net898),
    .X(_04306_));
 o211a_1 _18819_ (.A1(net740),
    .A2(_04306_),
    .B1(_04303_),
    .C1(net1497),
    .X(_04307_));
 a21oi_2 _18820_ (.A1(net68),
    .A2(net60),
    .B1(_04307_),
    .Y(_04308_));
 nand2_1 _18821_ (.A(net1471),
    .B(_04308_),
    .Y(_04309_));
 a32o_1 _18822_ (.A1(net1462),
    .A2(_04299_),
    .A3(_04309_),
    .B1(net1459),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[13] ),
    .X(_04310_));
 o22a_1 _18823_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[14] ),
    .A2(net1461),
    .B1(net1394),
    .B2(_04310_),
    .X(_00522_));
 mux2_1 _18824_ (.A0(\vmem_after_buf[63] ),
    .A1(\vmem_after_buf[47] ),
    .S(net925),
    .X(_04311_));
 mux2_1 _18825_ (.A0(\vmem_after_buf[31] ),
    .A1(\vmem_after_buf[15] ),
    .S(net925),
    .X(_04312_));
 mux2_1 _18826_ (.A0(_04311_),
    .A1(_04312_),
    .S(net908),
    .X(_04313_));
 mux2_1 _18827_ (.A0(\vmem_after_buf[95] ),
    .A1(\vmem_after_buf[79] ),
    .S(net925),
    .X(_04314_));
 mux2_1 _18828_ (.A0(\vmem_after_buf[127] ),
    .A1(\vmem_after_buf[111] ),
    .S(net925),
    .X(_04315_));
 mux2_1 _18829_ (.A0(_04314_),
    .A1(_04315_),
    .S(net894),
    .X(_04316_));
 mux2_1 _18830_ (.A0(_04313_),
    .A1(_04316_),
    .S(net731),
    .X(_04317_));
 mux2_1 _18831_ (.A0(net8),
    .A1(_04317_),
    .S(net1495),
    .X(_04318_));
 mux2_1 _18832_ (.A0(\vmem_after_buf[351] ),
    .A1(\vmem_after_buf[335] ),
    .S(net931),
    .X(_04319_));
 mux2_1 _18833_ (.A0(\vmem_after_buf[383] ),
    .A1(\vmem_after_buf[367] ),
    .S(net931),
    .X(_04320_));
 mux2_1 _18834_ (.A0(_04319_),
    .A1(_04320_),
    .S(net896),
    .X(_04321_));
 mux2_1 _18835_ (.A0(\vmem_after_buf[287] ),
    .A1(\vmem_after_buf[271] ),
    .S(net931),
    .X(_04322_));
 mux2_1 _18836_ (.A0(\vmem_after_buf[319] ),
    .A1(\vmem_after_buf[303] ),
    .S(net931),
    .X(_04323_));
 mux2_1 _18837_ (.A0(_04322_),
    .A1(_04323_),
    .S(net896),
    .X(_04324_));
 mux2_1 _18838_ (.A0(_04321_),
    .A1(_04324_),
    .S(net777),
    .X(_04325_));
 mux2_1 _18839_ (.A0(net43),
    .A1(_04325_),
    .S(net1497),
    .X(_04326_));
 mux2_1 _18840_ (.A0(\vmem_after_buf[223] ),
    .A1(\vmem_after_buf[207] ),
    .S(net926),
    .X(_04327_));
 mux2_1 _18841_ (.A0(\vmem_after_buf[255] ),
    .A1(\vmem_after_buf[239] ),
    .S(net925),
    .X(_04328_));
 mux2_1 _18842_ (.A0(_04327_),
    .A1(_04328_),
    .S(net893),
    .X(_04329_));
 mux2_1 _18843_ (.A0(\vmem_after_buf[159] ),
    .A1(\vmem_after_buf[143] ),
    .S(net925),
    .X(_04330_));
 mux2_1 _18844_ (.A0(\vmem_after_buf[191] ),
    .A1(\vmem_after_buf[175] ),
    .S(net926),
    .X(_04331_));
 mux2_1 _18845_ (.A0(_04330_),
    .A1(_04331_),
    .S(net894),
    .X(_04332_));
 mux2_1 _18846_ (.A0(_04329_),
    .A1(_04332_),
    .S(net773),
    .X(_04333_));
 mux2_1 _18847_ (.A0(net26),
    .A1(_04333_),
    .S(net1495),
    .X(_04334_));
 a22o_1 _18848_ (.A1(net1467),
    .A2(_04326_),
    .B1(_04334_),
    .B2(_03828_),
    .X(_04335_));
 a211o_1 _18849_ (.A1(net1468),
    .A2(_04318_),
    .B1(_04335_),
    .C1(net1471),
    .X(_04336_));
 or2_1 _18850_ (.A(\vmem_after_buf[463] ),
    .B(net953),
    .X(_04337_));
 o211a_1 _18851_ (.A1(\vmem_after_buf[479] ),
    .A2(net931),
    .B1(_04337_),
    .C1(net907),
    .X(_04338_));
 mux2_1 _18852_ (.A0(\vmem_after_buf[511] ),
    .A1(\vmem_after_buf[495] ),
    .S(net931),
    .X(_04339_));
 a211o_1 _18853_ (.A1(net896),
    .A2(_04339_),
    .B1(_04338_),
    .C1(net778),
    .X(_04340_));
 mux2_1 _18854_ (.A0(\vmem_after_buf[415] ),
    .A1(\vmem_after_buf[399] ),
    .S(net931),
    .X(_04341_));
 mux2_1 _18855_ (.A0(\vmem_after_buf[447] ),
    .A1(\vmem_after_buf[431] ),
    .S(net931),
    .X(_04342_));
 mux2_1 _18856_ (.A0(_04341_),
    .A1(_04342_),
    .S(net896),
    .X(_04343_));
 o211a_1 _18857_ (.A1(net736),
    .A2(_04343_),
    .B1(_04340_),
    .C1(net1497),
    .X(_04344_));
 a21oi_1 _18858_ (.A1(net68),
    .A2(net61),
    .B1(_04344_),
    .Y(_04345_));
 nand2_1 _18859_ (.A(net1471),
    .B(_04345_),
    .Y(_04346_));
 a32o_1 _18860_ (.A1(net1462),
    .A2(_04336_),
    .A3(_04346_),
    .B1(net1459),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[14] ),
    .X(_04347_));
 o22a_1 _18861_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[15] ),
    .A2(net1461),
    .B1(net1395),
    .B2(_04347_),
    .X(_00523_));
 or2_1 _18862_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[0] ),
    .B(_11017_),
    .X(_04348_));
 a21bo_1 _18863_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[0] ),
    .A2(_09644_),
    .B1_N(_04348_),
    .X(_00524_));
 xnor2_1 _18864_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[1] ),
    .B(_04348_),
    .Y(_00525_));
 or3_1 _18865_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[1] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[2] ),
    .C(_04348_),
    .X(_04349_));
 o21ai_1 _18866_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[1] ),
    .A2(_04348_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[2] ),
    .Y(_04350_));
 nand2_1 _18867_ (.A(_04349_),
    .B(_04350_),
    .Y(_00526_));
 xnor2_1 _18868_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[3] ),
    .B(_04349_),
    .Y(_00527_));
 o21a_1 _18869_ (.A1(_09642_),
    .A2(_04348_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[4] ),
    .X(_00528_));
 o21ai_1 _18870_ (.A1(_00113_),
    .A2(_10771_),
    .B1(_03752_),
    .Y(_04351_));
 nand2_1 _18871_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[0] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[1] ),
    .Y(_04352_));
 mux2_1 _18872_ (.A0(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[0] ),
    .A1(_04352_),
    .S(_04351_),
    .X(_00529_));
 nor3_1 _18873_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[0] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[1] ),
    .C(_03752_),
    .Y(_04353_));
 o21a_1 _18874_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[0] ),
    .A2(_03752_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[1] ),
    .X(_04354_));
 or3_1 _18875_ (.A(_10772_),
    .B(_04353_),
    .C(_04354_),
    .X(_00530_));
 or4_1 _18876_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[0] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[1] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[2] ),
    .D(_03752_),
    .X(_04355_));
 nand2b_1 _18877_ (.A_N(_04353_),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[2] ),
    .Y(_04356_));
 nand3b_1 _18878_ (.A_N(_10772_),
    .B(_04355_),
    .C(_04356_),
    .Y(_00531_));
 a21o_1 _18879_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[3] ),
    .A2(_04355_),
    .B1(_10772_),
    .X(_00532_));
 and2b_1 _18880_ (.A_N(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.mbist_end ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.form_end ),
    .X(_04357_));
 nor2_1 _18881_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.form_end ),
    .B(_09626_),
    .Y(_04358_));
 a221o_1 _18882_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[0] ),
    .A2(_04357_),
    .B1(_04358_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[0] ),
    .C1(net1464),
    .X(_04359_));
 o21a_1 _18883_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[0] ),
    .A2(_09631_),
    .B1(_04359_),
    .X(_00533_));
 a221o_1 _18884_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[1] ),
    .A2(_04357_),
    .B1(_04358_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[1] ),
    .C1(net1464),
    .X(_04360_));
 o21a_1 _18885_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[1] ),
    .A2(_09631_),
    .B1(_04360_),
    .X(_00534_));
 a221o_1 _18886_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[2] ),
    .A2(_04357_),
    .B1(_04358_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[2] ),
    .C1(net1464),
    .X(_04361_));
 o21a_1 _18887_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[2] ),
    .A2(_09631_),
    .B1(_04361_),
    .X(_00535_));
 a221o_1 _18888_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[3] ),
    .A2(_04357_),
    .B1(_04358_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[3] ),
    .C1(net1464),
    .X(_04362_));
 o21a_1 _18889_ (.A1(net1479),
    .A2(_09631_),
    .B1(_04362_),
    .X(_00536_));
 a221o_1 _18890_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[4] ),
    .A2(_04357_),
    .B1(_04358_),
    .B2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[4] ),
    .C1(net1464),
    .X(_04363_));
 o21a_1 _18891_ (.A1(net1477),
    .A2(_09631_),
    .B1(_04363_),
    .X(_00537_));
 or3_1 _18892_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[1] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[8] ),
    .C(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.mbist_end ),
    .X(_00538_));
 o21ba_1 _18893_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[8] ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.mbist_result ),
    .B1_N(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[1] ),
    .X(_00539_));
 mux2_1 _18894_ (.A0(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.read_after_prog_ok ),
    .A1(_09609_),
    .S(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_int_wr_bit ),
    .X(_00540_));
 nor2_1 _18895_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[8] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[6] ),
    .Y(_04364_));
 or2_1 _18896_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[0] ),
    .B(_04364_),
    .X(_04365_));
 nand2_1 _18897_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[0] ),
    .B(_04364_),
    .Y(_04366_));
 nand2_1 _18898_ (.A(_04365_),
    .B(_04366_),
    .Y(_00541_));
 xnor2_1 _18899_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[1] ),
    .B(_04365_),
    .Y(_00542_));
 or3_2 _18900_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[1] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[2] ),
    .C(_04365_),
    .X(_04367_));
 o21ai_1 _18901_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[1] ),
    .A2(_04365_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[2] ),
    .Y(_04368_));
 nand2_1 _18902_ (.A(_04367_),
    .B(_04368_),
    .Y(_00543_));
 xnor2_1 _18903_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[3] ),
    .B(_04367_),
    .Y(_00544_));
 or3_1 _18904_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[3] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[4] ),
    .C(_04367_),
    .X(_04369_));
 o21ai_1 _18905_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[3] ),
    .A2(_04367_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[4] ),
    .Y(_04370_));
 nand2_1 _18906_ (.A(_04369_),
    .B(_04370_),
    .Y(_00545_));
 or2_1 _18907_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[5] ),
    .B(_04369_),
    .X(_04371_));
 nand2_1 _18908_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[5] ),
    .B(_04369_),
    .Y(_04372_));
 nand2_1 _18909_ (.A(_04371_),
    .B(_04372_),
    .Y(_00546_));
 or2_1 _18910_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[6] ),
    .B(_04371_),
    .X(_04373_));
 nand2_1 _18911_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[6] ),
    .B(_04371_),
    .Y(_04374_));
 nand2_1 _18912_ (.A(_04373_),
    .B(_04374_),
    .Y(_00547_));
 or3_1 _18913_ (.A(_09617_),
    .B(_09618_),
    .C(_04364_),
    .X(_04375_));
 a21bo_1 _18914_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[7] ),
    .A2(_04373_),
    .B1_N(_04375_),
    .X(_00548_));
 xnor2_1 _18915_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[8] ),
    .B(_04375_),
    .Y(_00549_));
 o21a_1 _18916_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[8] ),
    .A2(_04375_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[9] ),
    .X(_04376_));
 a211o_1 _18917_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[8] ),
    .A2(_09619_),
    .B1(_09646_),
    .C1(_04376_),
    .X(_00550_));
 nor2_1 _18918_ (.A(net1502),
    .B(net1504),
    .Y(_04377_));
 o21bai_1 _18919_ (.A1(net1322),
    .A2(_04377_),
    .B1_N(\digitop_pav2.testctrl_pav2.inst_enter.tm_enter ),
    .Y(_00551_));
 o31ai_2 _18920_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[2] ),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[3] ),
    .A3(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[1] ),
    .B1(_09626_),
    .Y(_04378_));
 nand2_1 _18921_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[0] ),
    .B(_04378_),
    .Y(_04379_));
 or2_1 _18922_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[0] ),
    .B(_04378_),
    .X(_04380_));
 o21ai_1 _18923_ (.A1(_07159_),
    .A2(_04380_),
    .B1(_04379_),
    .Y(_00552_));
 or2_1 _18924_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[1] ),
    .B(_04380_),
    .X(_04381_));
 nand2_1 _18925_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[1] ),
    .B(_04380_),
    .Y(_04382_));
 nor2_2 _18926_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.reg_wr_en ),
    .B(_04378_),
    .Y(_04383_));
 a21oi_1 _18927_ (.A1(_04381_),
    .A2(_04382_),
    .B1(_04383_),
    .Y(_00553_));
 o21a_1 _18928_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[1] ),
    .A2(_04380_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[2] ),
    .X(_04384_));
 or3_1 _18929_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[1] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[2] ),
    .C(_04380_),
    .X(_04385_));
 or3b_1 _18930_ (.A(_04383_),
    .B(_04384_),
    .C_N(_04385_),
    .X(_00554_));
 or2_1 _18931_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[3] ),
    .B(_04385_),
    .X(_04386_));
 nand2_1 _18932_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[3] ),
    .B(_04385_),
    .Y(_04387_));
 a21oi_1 _18933_ (.A1(_04386_),
    .A2(_04387_),
    .B1(_04383_),
    .Y(_00555_));
 or3_1 _18934_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[3] ),
    .B(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[4] ),
    .C(_04385_),
    .X(_04388_));
 o21ai_1 _18935_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[3] ),
    .A2(_04385_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[4] ),
    .Y(_04389_));
 a21oi_1 _18936_ (.A1(_04388_),
    .A2(_04389_),
    .B1(_04383_),
    .Y(_00556_));
 or2_1 _18937_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[5] ),
    .B(_04388_),
    .X(_04390_));
 nand2_1 _18938_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[5] ),
    .B(_04388_),
    .Y(_04391_));
 a21oi_1 _18939_ (.A1(_04390_),
    .A2(_04391_),
    .B1(_04383_),
    .Y(_00557_));
 or2_1 _18940_ (.A(_09625_),
    .B(_04378_),
    .X(_04392_));
 nand2_1 _18941_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[6] ),
    .B(_04390_),
    .Y(_04393_));
 a21oi_1 _18942_ (.A1(_04392_),
    .A2(_04393_),
    .B1(_04383_),
    .Y(_00558_));
 or2_1 _18943_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[7] ),
    .B(_04392_),
    .X(_04394_));
 a21oi_1 _18944_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[7] ),
    .A2(_04392_),
    .B1(_04383_),
    .Y(_04395_));
 nand2_1 _18945_ (.A(_04394_),
    .B(_04395_),
    .Y(_00559_));
 or2_1 _18946_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[8] ),
    .B(_04394_),
    .X(_04396_));
 a21oi_1 _18947_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[8] ),
    .A2(_04394_),
    .B1(_04383_),
    .Y(_04397_));
 nand2_1 _18948_ (.A(_04396_),
    .B(_04397_),
    .Y(_00560_));
 a21o_1 _18949_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[9] ),
    .A2(_04396_),
    .B1(_04383_),
    .X(_00561_));
 a21o_1 _18950_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[3] ),
    .A2(_09609_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[2] ),
    .X(_04398_));
 a41o_1 _18951_ (.A1(net1480),
    .A2(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[4] ),
    .A3(_09592_),
    .A4(_09609_),
    .B1(_11012_),
    .X(_04399_));
 a31oi_1 _18952_ (.A1(net1480),
    .A2(_09612_),
    .A3(_04398_),
    .B1(_04399_),
    .Y(_04400_));
 or2_2 _18953_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[0] ),
    .B(_04400_),
    .X(_04401_));
 nand2_1 _18954_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[0] ),
    .B(_04400_),
    .Y(_04402_));
 nand2_1 _18955_ (.A(_04401_),
    .B(_04402_),
    .Y(_00562_));
 xnor2_1 _18956_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[1] ),
    .B(_04401_),
    .Y(_00563_));
 o21ai_1 _18957_ (.A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[1] ),
    .A2(_04401_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[2] ),
    .Y(_04403_));
 o21ai_1 _18958_ (.A1(_09590_),
    .A2(_04401_),
    .B1(_04403_),
    .Y(_00564_));
 or3_1 _18959_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[3] ),
    .B(_09590_),
    .C(_04401_),
    .X(_04404_));
 o21ai_1 _18960_ (.A1(_09590_),
    .A2(_04401_),
    .B1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[3] ),
    .Y(_04405_));
 nand2_1 _18961_ (.A(_04404_),
    .B(_04405_),
    .Y(_00565_));
 nand2_1 _18962_ (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[4] ),
    .B(_04404_),
    .Y(_04406_));
 o21ai_1 _18963_ (.A1(_09592_),
    .A2(_04400_),
    .B1(_04406_),
    .Y(_00566_));
 nand2_1 _18964_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[0] ),
    .B(_00161_),
    .Y(_00567_));
 nand2_1 _18965_ (.A(_11101_),
    .B(_00161_),
    .Y(_04407_));
 o21a_1 _18966_ (.A1(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[1] ),
    .A2(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[0] ),
    .B1(_04407_),
    .X(_00568_));
 mux2_1 _18967_ (.A0(_11101_),
    .A1(_04407_),
    .S(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[2] ),
    .X(_00569_));
 a31o_1 _18968_ (.A1(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[1] ),
    .A2(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[0] ),
    .A3(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[2] ),
    .B1(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[3] ),
    .X(_04408_));
 a21boi_1 _18969_ (.A1(_11102_),
    .A2(_00161_),
    .B1_N(_04408_),
    .Y(_00570_));
 nand2b_1 _18970_ (.A_N(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[5] ),
    .B(_11103_),
    .Y(_04409_));
 o21a_1 _18971_ (.A1(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[4] ),
    .A2(_11102_),
    .B1(_04409_),
    .X(_00571_));
 or2_1 _18972_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[5] ),
    .B(_11103_),
    .X(_00572_));
 o31ai_1 _18973_ (.A1(_07236_),
    .A2(\digitop_pav2.sync_inst.inst_rstx.gray_counter[0] ),
    .A3(\digitop_pav2.sync_inst.inst_rstx.gray_counter[1] ),
    .B1(net1400),
    .Y(_00573_));
 nor2_1 _18974_ (.A(net1399),
    .B(net1728),
    .Y(_00204_));
 nor2_1 _18975_ (.A(net1398),
    .B(net1250),
    .Y(_00214_));
 a21oi_1 _18976_ (.A1(net1247),
    .A2(\digitop_pav2.proc_ctrl_inst.cmdfsm.mode ),
    .B1(net1398),
    .Y(_00205_));
 nor2_1 _18977_ (.A(net1400),
    .B(net1832),
    .Y(_00208_));
 a21bo_1 _18978_ (.A1(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div4_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .A2(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_en.slow_clk_en_b_ff2_i ),
    .B1_N(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_en.slow_clk_en_b_ff3 ),
    .X(_04410_));
 o21a_1 _18979_ (.A1(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div4_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .A2(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_en.slow_clk_en_b_ff2_i ),
    .B1(_04410_),
    .X(_00578_));
 or2_1 _18980_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.en_scwend_clk_b ),
    .B(_11104_),
    .X(_00579_));
 a21o_1 _18981_ (.A1(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.en_pup_clk_b_aux ),
    .A2(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.en_pup_clk_b ),
    .B1(_11104_),
    .X(_00581_));
 and3_1 _18982_ (.A(net1456),
    .B(net1245),
    .C(_09160_),
    .X(_00213_));
 and2_1 _18983_ (.A(\digitop_pav2.sec_inst.ld_mem.st[0] ),
    .B(net1636),
    .X(_04411_));
 nand2_1 _18984_ (.A(\digitop_pav2.sec_inst.ld_mem.st[0] ),
    .B(net1636),
    .Y(_04412_));
 or3b_1 _18985_ (.A(\digitop_pav2.sec_inst.ld_mem.st[1] ),
    .B(_04411_),
    .C_N(\digitop_pav2.sec_inst.ld_mem.wctr[0] ),
    .X(_04413_));
 o21ai_1 _18986_ (.A1(\digitop_pav2.sec_inst.ld_mem.wctr[0] ),
    .A2(_04412_),
    .B1(_04413_),
    .Y(_00583_));
 nand2_1 _18987_ (.A(\digitop_pav2.sec_inst.ld_mem.wctr[0] ),
    .B(\digitop_pav2.sec_inst.ld_mem.wctr[1] ),
    .Y(_04414_));
 and3b_1 _18988_ (.A_N(\digitop_pav2.sec_inst.ld_mem.st[1] ),
    .B(_04412_),
    .C(\digitop_pav2.sec_inst.ld_mem.wctr[1] ),
    .X(_04415_));
 a31o_1 _18989_ (.A1(_09656_),
    .A2(_04411_),
    .A3(_04414_),
    .B1(_04415_),
    .X(_00584_));
 nor2_1 _18990_ (.A(_04412_),
    .B(_04414_),
    .Y(_04416_));
 and2_1 _18991_ (.A(\digitop_pav2.sec_inst.ld_mem.wctr[2] ),
    .B(_04416_),
    .X(_04417_));
 nor2_1 _18992_ (.A(\digitop_pav2.sec_inst.ld_mem.st[1] ),
    .B(_04417_),
    .Y(_04418_));
 o21a_1 _18993_ (.A1(\digitop_pav2.sec_inst.ld_mem.wctr[2] ),
    .A2(_04416_),
    .B1(_04418_),
    .X(_00585_));
 mux2_1 _18994_ (.A0(_04417_),
    .A1(_04418_),
    .S(\digitop_pav2.sec_inst.ld_mem.wctr[3] ),
    .X(_00586_));
 or4_1 _18995_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[6] ),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[11] ),
    .C(\digitop_pav2.rng_inst.rng_prngx_pav2.rngx_sec_req_i ),
    .D(\digitop_pav2.func_rnclk_en ),
    .X(_04419_));
 mux2_1 _18996_ (.A0(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[0] ),
    .A1(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[1] ),
    .S(net679),
    .X(_00587_));
 mux2_1 _18997_ (.A0(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[1] ),
    .A1(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[2] ),
    .S(net679),
    .X(_00588_));
 nand2_1 _18998_ (.A(\digitop_pav2.func_rnclk_en ),
    .B(\digitop_pav2.rng_inst.rng_prngx_pav2.trngx_data_i ),
    .Y(_04420_));
 xnor2_1 _18999_ (.A(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[0] ),
    .B(_04420_),
    .Y(_04421_));
 mux2_1 _19000_ (.A0(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[2] ),
    .A1(_04421_),
    .S(net679),
    .X(_00589_));
 a21oi_1 _19001_ (.A1(\digitop_pav2.sec_inst.ld_r.st[0] ),
    .A2(\digitop_pav2.sec_inst.ld_r.st[1] ),
    .B1(net716),
    .Y(_04422_));
 nor2_1 _19002_ (.A(_11412_),
    .B(_04422_),
    .Y(_00590_));
 and2_1 _19003_ (.A(_11405_),
    .B(_11413_),
    .X(_00591_));
 nand2_2 _19004_ (.A(\digitop_pav2.sec_inst.shift_in.st[2] ),
    .B(\digitop_pav2.sec_inst.shift_in.st[3] ),
    .Y(_04423_));
 nor2_1 _19005_ (.A(_03008_),
    .B(_04423_),
    .Y(_04424_));
 mux2_1 _19006_ (.A0(\digitop_pav2.sec_inst.reg160[16] ),
    .A1(net812),
    .S(net588),
    .X(_00592_));
 mux2_1 _19007_ (.A0(\digitop_pav2.sec_inst.reg160[17] ),
    .A1(\digitop_pav2.sec_inst.reg160[16] ),
    .S(net588),
    .X(_00593_));
 mux2_1 _19008_ (.A0(\digitop_pav2.sec_inst.reg160[18] ),
    .A1(\digitop_pav2.sec_inst.reg160[17] ),
    .S(net588),
    .X(_00594_));
 mux2_1 _19009_ (.A0(\digitop_pav2.sec_inst.reg160[19] ),
    .A1(\digitop_pav2.sec_inst.reg160[18] ),
    .S(net588),
    .X(_00595_));
 mux2_1 _19010_ (.A0(\digitop_pav2.sec_inst.reg160[20] ),
    .A1(\digitop_pav2.sec_inst.reg160[19] ),
    .S(net588),
    .X(_00596_));
 mux2_1 _19011_ (.A0(\digitop_pav2.sec_inst.reg160[21] ),
    .A1(\digitop_pav2.sec_inst.reg160[20] ),
    .S(net588),
    .X(_00597_));
 mux2_1 _19012_ (.A0(\digitop_pav2.sec_inst.reg160[22] ),
    .A1(\digitop_pav2.sec_inst.reg160[21] ),
    .S(net588),
    .X(_00598_));
 mux2_1 _19013_ (.A0(\digitop_pav2.sec_inst.reg160[23] ),
    .A1(\digitop_pav2.sec_inst.reg160[22] ),
    .S(net589),
    .X(_00599_));
 mux2_1 _19014_ (.A0(\digitop_pav2.sec_inst.reg160[24] ),
    .A1(\digitop_pav2.sec_inst.reg160[23] ),
    .S(net588),
    .X(_00600_));
 mux2_1 _19015_ (.A0(\digitop_pav2.sec_inst.reg160[25] ),
    .A1(\digitop_pav2.sec_inst.reg160[24] ),
    .S(net588),
    .X(_00601_));
 mux2_1 _19016_ (.A0(\digitop_pav2.sec_inst.reg160[26] ),
    .A1(\digitop_pav2.sec_inst.reg160[25] ),
    .S(net589),
    .X(_00602_));
 mux2_1 _19017_ (.A0(\digitop_pav2.sec_inst.reg160[27] ),
    .A1(\digitop_pav2.sec_inst.reg160[26] ),
    .S(net589),
    .X(_00603_));
 mux2_1 _19018_ (.A0(\digitop_pav2.sec_inst.reg160[28] ),
    .A1(\digitop_pav2.sec_inst.reg160[27] ),
    .S(net589),
    .X(_00604_));
 mux2_1 _19019_ (.A0(\digitop_pav2.sec_inst.reg160[29] ),
    .A1(\digitop_pav2.sec_inst.reg160[28] ),
    .S(net589),
    .X(_00605_));
 mux2_1 _19020_ (.A0(\digitop_pav2.sec_inst.reg160[30] ),
    .A1(\digitop_pav2.sec_inst.reg160[29] ),
    .S(net589),
    .X(_00606_));
 mux2_1 _19021_ (.A0(\digitop_pav2.sec_inst.reg160[31] ),
    .A1(\digitop_pav2.sec_inst.reg160[30] ),
    .S(net589),
    .X(_00607_));
 nor2_1 _19022_ (.A(_11409_),
    .B(_04423_),
    .Y(_04425_));
 mux2_1 _19023_ (.A0(\digitop_pav2.sec_inst.reg160[32] ),
    .A1(net812),
    .S(net586),
    .X(_00608_));
 mux2_1 _19024_ (.A0(\digitop_pav2.sec_inst.reg160[33] ),
    .A1(\digitop_pav2.sec_inst.reg160[32] ),
    .S(net586),
    .X(_00609_));
 mux2_1 _19025_ (.A0(\digitop_pav2.sec_inst.reg160[34] ),
    .A1(\digitop_pav2.sec_inst.reg160[33] ),
    .S(net586),
    .X(_00610_));
 mux2_1 _19026_ (.A0(\digitop_pav2.sec_inst.reg160[35] ),
    .A1(\digitop_pav2.sec_inst.reg160[34] ),
    .S(net586),
    .X(_00611_));
 mux2_1 _19027_ (.A0(\digitop_pav2.sec_inst.reg160[36] ),
    .A1(\digitop_pav2.sec_inst.reg160[35] ),
    .S(net586),
    .X(_00612_));
 mux2_1 _19028_ (.A0(\digitop_pav2.sec_inst.reg160[37] ),
    .A1(\digitop_pav2.sec_inst.reg160[36] ),
    .S(net586),
    .X(_00613_));
 mux2_1 _19029_ (.A0(\digitop_pav2.sec_inst.reg160[38] ),
    .A1(\digitop_pav2.sec_inst.reg160[37] ),
    .S(net586),
    .X(_00614_));
 mux2_1 _19030_ (.A0(\digitop_pav2.sec_inst.reg160[39] ),
    .A1(\digitop_pav2.sec_inst.reg160[38] ),
    .S(net586),
    .X(_00615_));
 mux2_1 _19031_ (.A0(\digitop_pav2.sec_inst.reg160[40] ),
    .A1(\digitop_pav2.sec_inst.reg160[39] ),
    .S(net586),
    .X(_00616_));
 mux2_1 _19032_ (.A0(\digitop_pav2.sec_inst.reg160[41] ),
    .A1(\digitop_pav2.sec_inst.reg160[40] ),
    .S(net586),
    .X(_00617_));
 mux2_1 _19033_ (.A0(\digitop_pav2.sec_inst.reg160[42] ),
    .A1(\digitop_pav2.sec_inst.reg160[41] ),
    .S(net587),
    .X(_00618_));
 mux2_1 _19034_ (.A0(\digitop_pav2.sec_inst.reg160[43] ),
    .A1(\digitop_pav2.sec_inst.reg160[42] ),
    .S(net587),
    .X(_00619_));
 mux2_1 _19035_ (.A0(\digitop_pav2.sec_inst.reg160[44] ),
    .A1(\digitop_pav2.sec_inst.reg160[43] ),
    .S(net587),
    .X(_00620_));
 mux2_1 _19036_ (.A0(\digitop_pav2.sec_inst.reg160[45] ),
    .A1(\digitop_pav2.sec_inst.reg160[44] ),
    .S(net587),
    .X(_00621_));
 mux2_1 _19037_ (.A0(\digitop_pav2.sec_inst.reg160[46] ),
    .A1(\digitop_pav2.sec_inst.reg160[45] ),
    .S(net587),
    .X(_00622_));
 mux2_1 _19038_ (.A0(\digitop_pav2.sec_inst.reg160[47] ),
    .A1(\digitop_pav2.sec_inst.reg160[46] ),
    .S(net587),
    .X(_00623_));
 nor2_1 _19039_ (.A(_03004_),
    .B(_04423_),
    .Y(_04426_));
 mux2_1 _19040_ (.A0(\digitop_pav2.sec_inst.reg160[48] ),
    .A1(net812),
    .S(net585),
    .X(_00624_));
 mux2_1 _19041_ (.A0(\digitop_pav2.sec_inst.reg160[49] ),
    .A1(\digitop_pav2.sec_inst.reg160[48] ),
    .S(net585),
    .X(_00625_));
 mux2_1 _19042_ (.A0(\digitop_pav2.sec_inst.reg160[50] ),
    .A1(\digitop_pav2.sec_inst.reg160[49] ),
    .S(net584),
    .X(_00626_));
 mux2_1 _19043_ (.A0(\digitop_pav2.sec_inst.reg160[51] ),
    .A1(\digitop_pav2.sec_inst.reg160[50] ),
    .S(net584),
    .X(_00627_));
 mux2_1 _19044_ (.A0(\digitop_pav2.sec_inst.reg160[52] ),
    .A1(\digitop_pav2.sec_inst.reg160[51] ),
    .S(net584),
    .X(_00628_));
 mux2_1 _19045_ (.A0(\digitop_pav2.sec_inst.reg160[53] ),
    .A1(\digitop_pav2.sec_inst.reg160[52] ),
    .S(net584),
    .X(_00629_));
 mux2_1 _19046_ (.A0(\digitop_pav2.sec_inst.reg160[54] ),
    .A1(\digitop_pav2.sec_inst.reg160[53] ),
    .S(net585),
    .X(_00630_));
 mux2_1 _19047_ (.A0(\digitop_pav2.sec_inst.reg160[55] ),
    .A1(\digitop_pav2.sec_inst.reg160[54] ),
    .S(net584),
    .X(_00631_));
 mux2_1 _19048_ (.A0(\digitop_pav2.sec_inst.reg160[56] ),
    .A1(\digitop_pav2.sec_inst.reg160[55] ),
    .S(net584),
    .X(_00632_));
 mux2_1 _19049_ (.A0(\digitop_pav2.sec_inst.reg160[57] ),
    .A1(\digitop_pav2.sec_inst.reg160[56] ),
    .S(net584),
    .X(_00633_));
 mux2_1 _19050_ (.A0(\digitop_pav2.sec_inst.reg160[58] ),
    .A1(\digitop_pav2.sec_inst.reg160[57] ),
    .S(net585),
    .X(_00634_));
 mux2_1 _19051_ (.A0(\digitop_pav2.sec_inst.reg160[59] ),
    .A1(\digitop_pav2.sec_inst.reg160[58] ),
    .S(net585),
    .X(_00635_));
 mux2_1 _19052_ (.A0(\digitop_pav2.sec_inst.reg160[60] ),
    .A1(\digitop_pav2.sec_inst.reg160[59] ),
    .S(net584),
    .X(_00636_));
 mux2_1 _19053_ (.A0(\digitop_pav2.sec_inst.reg160[61] ),
    .A1(\digitop_pav2.sec_inst.reg160[60] ),
    .S(net584),
    .X(_00637_));
 mux2_1 _19054_ (.A0(\digitop_pav2.sec_inst.reg160[62] ),
    .A1(\digitop_pav2.sec_inst.reg160[61] ),
    .S(net584),
    .X(_00638_));
 mux2_1 _19055_ (.A0(\digitop_pav2.sec_inst.reg160[63] ),
    .A1(\digitop_pav2.sec_inst.reg160[62] ),
    .S(net585),
    .X(_00639_));
 mux2_1 _19056_ (.A0(\digitop_pav2.sec_inst.shift_in.s12.q[0] ),
    .A1(net1641),
    .S(_11425_),
    .X(_00640_));
 mux2_1 _19057_ (.A0(\digitop_pav2.sec_inst.shift_in.s12.q[0] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s12.q[1] ),
    .S(_11424_),
    .X(_00641_));
 mux2_1 _19058_ (.A0(\digitop_pav2.sec_inst.shift_in.s12.q[1] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s12.q[2] ),
    .S(_11424_),
    .X(_00642_));
 mux2_1 _19059_ (.A0(\digitop_pav2.sec_inst.shift_in.s12.q[2] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s12.q[3] ),
    .S(_11424_),
    .X(_00643_));
 mux2_1 _19060_ (.A0(\digitop_pav2.sec_inst.shift_in.s12.q[3] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s12.q[4] ),
    .S(_11424_),
    .X(_00644_));
 mux2_1 _19061_ (.A0(\digitop_pav2.sec_inst.shift_in.s12.q[4] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s12.q[5] ),
    .S(_11424_),
    .X(_00645_));
 mux2_1 _19062_ (.A0(\digitop_pav2.sec_inst.shift_in.s12.q[5] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[6] ),
    .S(_11424_),
    .X(_00646_));
 mux2_1 _19063_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[6] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[7] ),
    .S(_11424_),
    .X(_00647_));
 mux2_1 _19064_ (.A0(\digitop_pav2.sec_inst.shift_in.s11.q[0] ),
    .A1(net1641),
    .S(_03020_),
    .X(_00648_));
 mux2_1 _19065_ (.A0(\digitop_pav2.sec_inst.shift_in.s11.q[0] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s11.q[1] ),
    .S(_03021_),
    .X(_00649_));
 mux2_1 _19066_ (.A0(\digitop_pav2.sec_inst.shift_in.s11.q[1] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s11.q[2] ),
    .S(_03021_),
    .X(_00650_));
 mux2_1 _19067_ (.A0(\digitop_pav2.sec_inst.shift_in.s11.q[2] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s11.q[3] ),
    .S(_03021_),
    .X(_00651_));
 mux2_1 _19068_ (.A0(\digitop_pav2.sec_inst.shift_in.s11.q[3] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s11.q[4] ),
    .S(_03021_),
    .X(_00652_));
 mux2_1 _19069_ (.A0(\digitop_pav2.sec_inst.shift_in.s11.q[4] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s11.q[5] ),
    .S(_03021_),
    .X(_00653_));
 mux2_1 _19070_ (.A0(\digitop_pav2.sec_inst.shift_in.s11.q[5] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[14] ),
    .S(_03021_),
    .X(_00654_));
 mux2_1 _19071_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[15] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[14] ),
    .S(_03020_),
    .X(_00655_));
 mux2_1 _19072_ (.A0(\digitop_pav2.sec_inst.shift_in.s10.q[0] ),
    .A1(net812),
    .S(_11427_),
    .X(_00656_));
 mux2_1 _19073_ (.A0(\digitop_pav2.sec_inst.shift_in.s10.q[1] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s10.q[0] ),
    .S(_11427_),
    .X(_00657_));
 mux2_1 _19074_ (.A0(\digitop_pav2.sec_inst.shift_in.s10.q[2] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s10.q[1] ),
    .S(_11427_),
    .X(_00658_));
 mux2_1 _19075_ (.A0(\digitop_pav2.sec_inst.shift_in.s10.q[3] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s10.q[2] ),
    .S(_11427_),
    .X(_00659_));
 mux2_1 _19076_ (.A0(\digitop_pav2.sec_inst.shift_in.s10.q[4] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s10.q[3] ),
    .S(_11427_),
    .X(_00660_));
 mux2_1 _19077_ (.A0(\digitop_pav2.sec_inst.shift_in.s10.q[5] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s10.q[4] ),
    .S(_11427_),
    .X(_00661_));
 mux2_1 _19078_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[22] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s10.q[5] ),
    .S(_11427_),
    .X(_00662_));
 mux2_1 _19079_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[23] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[22] ),
    .S(_11427_),
    .X(_00663_));
 mux2_1 _19080_ (.A0(\digitop_pav2.sec_inst.shift_in.s1.q[0] ),
    .A1(net812),
    .S(_03005_),
    .X(_00664_));
 mux2_1 _19081_ (.A0(\digitop_pav2.sec_inst.shift_in.s1.q[0] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s1.q[1] ),
    .S(net593),
    .X(_00665_));
 mux2_1 _19082_ (.A0(\digitop_pav2.sec_inst.shift_in.s1.q[1] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s1.q[2] ),
    .S(net593),
    .X(_00666_));
 mux2_1 _19083_ (.A0(\digitop_pav2.sec_inst.shift_in.s1.q[2] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s1.q[3] ),
    .S(net593),
    .X(_00667_));
 mux2_1 _19084_ (.A0(\digitop_pav2.sec_inst.shift_in.s1.q[3] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s1.q[4] ),
    .S(net593),
    .X(_00668_));
 mux2_1 _19085_ (.A0(\digitop_pav2.sec_inst.shift_in.s1.q[4] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s1.q[5] ),
    .S(net593),
    .X(_00669_));
 mux2_1 _19086_ (.A0(\digitop_pav2.sec_inst.shift_in.s1.q[5] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[94] ),
    .S(net593),
    .X(_00670_));
 mux2_1 _19087_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[95] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[94] ),
    .S(_03005_),
    .X(_00671_));
 mux2_1 _19088_ (.A0(\digitop_pav2.sec_inst.shift_in.s8.q[0] ),
    .A1(net1641),
    .S(_11435_),
    .X(_00672_));
 mux2_1 _19089_ (.A0(\digitop_pav2.sec_inst.shift_in.s8.q[0] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s8.q[1] ),
    .S(net574),
    .X(_00673_));
 mux2_1 _19090_ (.A0(\digitop_pav2.sec_inst.shift_in.s8.q[1] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s8.q[2] ),
    .S(_11434_),
    .X(_00674_));
 mux2_1 _19091_ (.A0(\digitop_pav2.sec_inst.shift_in.s8.q[2] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s8.q[3] ),
    .S(_11434_),
    .X(_00675_));
 mux2_1 _19092_ (.A0(\digitop_pav2.sec_inst.shift_in.s8.q[3] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s8.q[4] ),
    .S(_11434_),
    .X(_00676_));
 mux2_1 _19093_ (.A0(\digitop_pav2.sec_inst.shift_in.s8.q[4] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s8.q[5] ),
    .S(_11434_),
    .X(_00677_));
 mux2_1 _19094_ (.A0(\digitop_pav2.sec_inst.shift_in.s8.q[5] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[38] ),
    .S(net574),
    .X(_00678_));
 mux2_1 _19095_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[38] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[39] ),
    .S(net574),
    .X(_00679_));
 a21bo_1 _19096_ (.A1(net1641),
    .A2(_03015_),
    .B1_N(_03016_),
    .X(_00680_));
 mux2_1 _19097_ (.A0(\digitop_pav2.sec_inst.shift_in.s7.q[1] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s7.q[0] ),
    .S(_03015_),
    .X(_00681_));
 mux2_1 _19098_ (.A0(\digitop_pav2.sec_inst.shift_in.s7.q[2] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s7.q[1] ),
    .S(_03015_),
    .X(_00682_));
 mux2_1 _19099_ (.A0(\digitop_pav2.sec_inst.shift_in.s7.q[3] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s7.q[2] ),
    .S(_03015_),
    .X(_00683_));
 mux2_1 _19100_ (.A0(\digitop_pav2.sec_inst.shift_in.s7.q[4] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s7.q[3] ),
    .S(_03015_),
    .X(_00684_));
 mux2_1 _19101_ (.A0(\digitop_pav2.sec_inst.shift_in.s7.q[5] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s7.q[4] ),
    .S(_03015_),
    .X(_00685_));
 mux2_1 _19102_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[46] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s7.q[5] ),
    .S(_03015_),
    .X(_00686_));
 mux2_1 _19103_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[47] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[46] ),
    .S(_03015_),
    .X(_00687_));
 mux2_1 _19104_ (.A0(\digitop_pav2.sec_inst.shift_in.s6.q[0] ),
    .A1(net812),
    .S(_11419_),
    .X(_00688_));
 mux2_1 _19105_ (.A0(\digitop_pav2.sec_inst.shift_in.s6.q[0] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s6.q[1] ),
    .S(net594),
    .X(_00689_));
 mux2_1 _19106_ (.A0(\digitop_pav2.sec_inst.shift_in.s6.q[1] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s6.q[2] ),
    .S(net594),
    .X(_00690_));
 mux2_1 _19107_ (.A0(\digitop_pav2.sec_inst.shift_in.s6.q[2] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s6.q[3] ),
    .S(net594),
    .X(_00691_));
 mux2_1 _19108_ (.A0(\digitop_pav2.sec_inst.shift_in.s6.q[3] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s6.q[4] ),
    .S(net594),
    .X(_00692_));
 mux2_1 _19109_ (.A0(\digitop_pav2.sec_inst.shift_in.s6.q[4] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s6.q[5] ),
    .S(net594),
    .X(_00693_));
 mux2_1 _19110_ (.A0(\digitop_pav2.sec_inst.shift_in.s6.q[5] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[54] ),
    .S(_11420_),
    .X(_00694_));
 mux2_1 _19111_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[55] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[54] ),
    .S(_11419_),
    .X(_00695_));
 mux2_1 _19112_ (.A0(\digitop_pav2.sec_inst.shift_in.s5.q[0] ),
    .A1(net1641),
    .S(_03012_),
    .X(_00696_));
 mux2_1 _19113_ (.A0(\digitop_pav2.sec_inst.shift_in.s5.q[0] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s5.q[1] ),
    .S(net591),
    .X(_00697_));
 mux2_1 _19114_ (.A0(\digitop_pav2.sec_inst.shift_in.s5.q[1] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s5.q[2] ),
    .S(net591),
    .X(_00698_));
 mux2_1 _19115_ (.A0(\digitop_pav2.sec_inst.shift_in.s5.q[2] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s5.q[3] ),
    .S(net591),
    .X(_00699_));
 mux2_1 _19116_ (.A0(\digitop_pav2.sec_inst.shift_in.s5.q[3] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s5.q[4] ),
    .S(net591),
    .X(_00700_));
 mux2_1 _19117_ (.A0(\digitop_pav2.sec_inst.shift_in.s5.q[4] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s5.q[5] ),
    .S(net591),
    .X(_00701_));
 mux2_1 _19118_ (.A0(\digitop_pav2.sec_inst.shift_in.s5.q[5] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[62] ),
    .S(_03013_),
    .X(_00702_));
 mux2_1 _19119_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[63] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[62] ),
    .S(_03012_),
    .X(_00703_));
 mux2_1 _19120_ (.A0(\digitop_pav2.sec_inst.shift_in.s4.q[0] ),
    .A1(net812),
    .S(_11402_),
    .X(_00704_));
 mux2_1 _19121_ (.A0(\digitop_pav2.sec_inst.shift_in.s4.q[0] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s4.q[1] ),
    .S(net577),
    .X(_00705_));
 mux2_1 _19122_ (.A0(\digitop_pav2.sec_inst.shift_in.s4.q[1] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s4.q[2] ),
    .S(net577),
    .X(_00706_));
 mux2_1 _19123_ (.A0(\digitop_pav2.sec_inst.shift_in.s4.q[2] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s4.q[3] ),
    .S(net577),
    .X(_00707_));
 mux2_1 _19124_ (.A0(\digitop_pav2.sec_inst.shift_in.s4.q[3] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s4.q[4] ),
    .S(_11401_),
    .X(_00708_));
 mux2_1 _19125_ (.A0(\digitop_pav2.sec_inst.shift_in.s4.q[4] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s4.q[5] ),
    .S(net577),
    .X(_00709_));
 mux2_1 _19126_ (.A0(\digitop_pav2.sec_inst.shift_in.s4.q[5] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[70] ),
    .S(net577),
    .X(_00710_));
 mux2_1 _19127_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[70] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[71] ),
    .S(net577),
    .X(_00711_));
 mux2_1 _19128_ (.A0(\digitop_pav2.sec_inst.shift_in.s3.q[0] ),
    .A1(net812),
    .S(_03009_),
    .X(_00712_));
 mux2_1 _19129_ (.A0(\digitop_pav2.sec_inst.shift_in.s3.q[0] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s3.q[1] ),
    .S(_03010_),
    .X(_00713_));
 mux2_1 _19130_ (.A0(\digitop_pav2.sec_inst.shift_in.s3.q[1] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s3.q[2] ),
    .S(net592),
    .X(_00714_));
 mux2_1 _19131_ (.A0(\digitop_pav2.sec_inst.shift_in.s3.q[2] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s3.q[3] ),
    .S(net592),
    .X(_00715_));
 mux2_1 _19132_ (.A0(\digitop_pav2.sec_inst.shift_in.s3.q[3] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s3.q[4] ),
    .S(net592),
    .X(_00716_));
 mux2_1 _19133_ (.A0(\digitop_pav2.sec_inst.shift_in.s3.q[4] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s3.q[5] ),
    .S(net592),
    .X(_00717_));
 mux2_1 _19134_ (.A0(\digitop_pav2.sec_inst.shift_in.s3.q[5] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[78] ),
    .S(net592),
    .X(_00718_));
 mux2_1 _19135_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[79] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[78] ),
    .S(_03009_),
    .X(_00719_));
 mux2_1 _19136_ (.A0(\digitop_pav2.sec_inst.shift_in.s2.q[0] ),
    .A1(net812),
    .S(_11410_),
    .X(_00720_));
 mux2_1 _19137_ (.A0(\digitop_pav2.sec_inst.shift_in.s2.q[0] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s2.q[1] ),
    .S(_11411_),
    .X(_00721_));
 mux2_1 _19138_ (.A0(\digitop_pav2.sec_inst.shift_in.s2.q[1] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s2.q[2] ),
    .S(net599),
    .X(_00722_));
 mux2_1 _19139_ (.A0(\digitop_pav2.sec_inst.shift_in.s2.q[2] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s2.q[3] ),
    .S(net599),
    .X(_00723_));
 mux2_1 _19140_ (.A0(\digitop_pav2.sec_inst.shift_in.s2.q[3] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s2.q[4] ),
    .S(net599),
    .X(_00724_));
 mux2_1 _19141_ (.A0(\digitop_pav2.sec_inst.shift_in.s2.q[4] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s2.q[5] ),
    .S(net599),
    .X(_00725_));
 mux2_1 _19142_ (.A0(\digitop_pav2.sec_inst.shift_in.s2.q[5] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[86] ),
    .S(net599),
    .X(_00726_));
 mux2_1 _19143_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[87] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[86] ),
    .S(_11410_),
    .X(_00727_));
 or2_1 _19144_ (.A(_11399_),
    .B(_04423_),
    .X(_04427_));
 inv_2 _19145_ (.A(net573),
    .Y(_04428_));
 mux2_1 _19146_ (.A0(\digitop_pav2.sec_inst.reg160[0] ),
    .A1(net812),
    .S(_04428_),
    .X(_00728_));
 mux2_1 _19147_ (.A0(\digitop_pav2.sec_inst.reg160[0] ),
    .A1(\digitop_pav2.sec_inst.reg160[1] ),
    .S(net572),
    .X(_00729_));
 mux2_1 _19148_ (.A0(\digitop_pav2.sec_inst.reg160[1] ),
    .A1(\digitop_pav2.sec_inst.reg160[2] ),
    .S(net572),
    .X(_00730_));
 mux2_1 _19149_ (.A0(\digitop_pav2.sec_inst.reg160[2] ),
    .A1(\digitop_pav2.sec_inst.reg160[3] ),
    .S(net572),
    .X(_00731_));
 mux2_1 _19150_ (.A0(\digitop_pav2.sec_inst.reg160[3] ),
    .A1(\digitop_pav2.sec_inst.reg160[4] ),
    .S(net572),
    .X(_00732_));
 mux2_1 _19151_ (.A0(\digitop_pav2.sec_inst.reg160[4] ),
    .A1(\digitop_pav2.sec_inst.reg160[5] ),
    .S(net572),
    .X(_00733_));
 mux2_1 _19152_ (.A0(\digitop_pav2.sec_inst.reg160[5] ),
    .A1(\digitop_pav2.sec_inst.reg160[6] ),
    .S(net572),
    .X(_00734_));
 mux2_1 _19153_ (.A0(\digitop_pav2.sec_inst.reg160[6] ),
    .A1(\digitop_pav2.sec_inst.reg160[7] ),
    .S(net572),
    .X(_00735_));
 mux2_1 _19154_ (.A0(\digitop_pav2.sec_inst.reg160[7] ),
    .A1(\digitop_pav2.sec_inst.reg160[8] ),
    .S(net572),
    .X(_00736_));
 mux2_1 _19155_ (.A0(\digitop_pav2.sec_inst.reg160[8] ),
    .A1(\digitop_pav2.sec_inst.reg160[9] ),
    .S(net573),
    .X(_00737_));
 mux2_1 _19156_ (.A0(\digitop_pav2.sec_inst.reg160[9] ),
    .A1(\digitop_pav2.sec_inst.reg160[10] ),
    .S(net572),
    .X(_00738_));
 mux2_1 _19157_ (.A0(\digitop_pav2.sec_inst.reg160[10] ),
    .A1(\digitop_pav2.sec_inst.reg160[11] ),
    .S(net572),
    .X(_00739_));
 mux2_1 _19158_ (.A0(\digitop_pav2.sec_inst.reg160[11] ),
    .A1(\digitop_pav2.sec_inst.reg160[12] ),
    .S(net573),
    .X(_00740_));
 mux2_1 _19159_ (.A0(\digitop_pav2.sec_inst.reg160[12] ),
    .A1(\digitop_pav2.sec_inst.reg160[13] ),
    .S(net573),
    .X(_00741_));
 mux2_1 _19160_ (.A0(\digitop_pav2.sec_inst.reg160[13] ),
    .A1(\digitop_pav2.sec_inst.reg160[14] ),
    .S(net573),
    .X(_00742_));
 mux2_1 _19161_ (.A0(\digitop_pav2.sec_inst.reg160[14] ),
    .A1(\digitop_pav2.sec_inst.reg160[15] ),
    .S(net573),
    .X(_00743_));
 a22o_1 _19162_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[55] ),
    .A2(_11419_),
    .B1(_11435_),
    .B2(\digitop_pav2.sec_inst.ld_r.reg96_i[39] ),
    .X(_04429_));
 a22o_1 _19163_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[87] ),
    .A2(_11410_),
    .B1(net587),
    .B2(\digitop_pav2.sec_inst.reg160[47] ),
    .X(_04430_));
 a221o_1 _19164_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[7] ),
    .A2(_11425_),
    .B1(_03009_),
    .B2(\digitop_pav2.sec_inst.ld_r.reg96_i[79] ),
    .C1(_04429_),
    .X(_04431_));
 a22o_1 _19165_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[63] ),
    .A2(_03012_),
    .B1(net590),
    .B2(\digitop_pav2.sec_inst.ld_r.reg96_i[31] ),
    .X(_04432_));
 a221o_1 _19166_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[47] ),
    .A2(_03015_),
    .B1(_04428_),
    .B2(\digitop_pav2.sec_inst.reg160[15] ),
    .C1(_04432_),
    .X(_04433_));
 a221o_1 _19167_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[95] ),
    .A2(_03005_),
    .B1(net588),
    .B2(\digitop_pav2.sec_inst.reg160[31] ),
    .C1(_04430_),
    .X(_04434_));
 a22o_1 _19168_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[23] ),
    .A2(_11427_),
    .B1(net585),
    .B2(\digitop_pav2.sec_inst.reg160[63] ),
    .X(_04435_));
 a221o_1 _19169_ (.A1(\digitop_pav2.sec_inst.ld_r.reg96_i[71] ),
    .A2(_11402_),
    .B1(_03020_),
    .B2(\digitop_pav2.sec_inst.ld_r.reg96_i[15] ),
    .C1(_04435_),
    .X(_04436_));
 or3_1 _19170_ (.A(_04433_),
    .B(_04434_),
    .C(_04436_),
    .X(_04437_));
 nor3_2 _19171_ (.A(net1646),
    .B(_04431_),
    .C(_04437_),
    .Y(_04438_));
 inv_2 _19172_ (.A(_04438_),
    .Y(_04439_));
 nand2_1 _19173_ (.A(\digitop_pav2.sec_inst.shift_in.st[0] ),
    .B(_04439_),
    .Y(_04440_));
 a21o_1 _19174_ (.A1(_03700_),
    .A2(_04439_),
    .B1(\digitop_pav2.sec_inst.shift_in.st[0] ),
    .X(_04441_));
 and2_1 _19175_ (.A(_04440_),
    .B(_04441_),
    .X(_00744_));
 nor2_1 _19176_ (.A(\digitop_pav2.sec_inst.shift_in.st[1] ),
    .B(_04438_),
    .Y(_04442_));
 a22o_1 _19177_ (.A1(\digitop_pav2.sec_inst.shift_in.st[1] ),
    .A2(_04440_),
    .B1(_04442_),
    .B2(\digitop_pav2.sec_inst.shift_in.st[0] ),
    .X(_00745_));
 nor2_1 _19178_ (.A(_11398_),
    .B(_04438_),
    .Y(_04443_));
 xor2_1 _19179_ (.A(\digitop_pav2.sec_inst.shift_in.st[2] ),
    .B(_04443_),
    .X(_00746_));
 a21o_1 _19180_ (.A1(\digitop_pav2.sec_inst.shift_in.st[2] ),
    .A2(_04443_),
    .B1(\digitop_pav2.sec_inst.shift_in.st[3] ),
    .X(_04444_));
 o31a_1 _19181_ (.A1(_11398_),
    .A2(_04423_),
    .A3(_04438_),
    .B1(_04444_),
    .X(_00747_));
 o31a_1 _19182_ (.A1(_11398_),
    .A2(_04423_),
    .A3(_04438_),
    .B1(\digitop_pav2.sec_inst.shift_in.st[4] ),
    .X(_04445_));
 a21o_1 _19183_ (.A1(_04428_),
    .A2(_04439_),
    .B1(_04445_),
    .X(_00748_));
 nor2_1 _19184_ (.A(net697),
    .B(_07523_),
    .Y(_04446_));
 a22o_1 _19185_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[0] ),
    .A2(net696),
    .B1(net331),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[0] ),
    .X(_00749_));
 a22o_1 _19186_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[1] ),
    .A2(net696),
    .B1(net331),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[1] ),
    .X(_00750_));
 a22o_1 _19187_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[2] ),
    .A2(net698),
    .B1(net333),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ),
    .X(_00751_));
 a22o_1 _19188_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[3] ),
    .A2(net696),
    .B1(net331),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[3] ),
    .X(_00752_));
 a22o_1 _19189_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[4] ),
    .A2(net698),
    .B1(net333),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[4] ),
    .X(_00753_));
 a22o_1 _19190_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[5] ),
    .A2(net696),
    .B1(net331),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[5] ),
    .X(_00754_));
 a22o_1 _19191_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[6] ),
    .A2(net696),
    .B1(net331),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[6] ),
    .X(_00755_));
 mux2_1 _19192_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[7] ),
    .A1(_08331_),
    .S(net711),
    .X(_00756_));
 a22o_1 _19193_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[8] ),
    .A2(net692),
    .B1(net324),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[8] ),
    .X(_00757_));
 a22o_1 _19194_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[9] ),
    .A2(net690),
    .B1(net328),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[9] ),
    .X(_00758_));
 a22o_1 _19195_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[10] ),
    .A2(net688),
    .B1(net324),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[10] ),
    .X(_00759_));
 a22o_1 _19196_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[11] ),
    .A2(net690),
    .B1(net327),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[11] ),
    .X(_00760_));
 a22o_1 _19197_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[12] ),
    .A2(net690),
    .B1(net327),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[12] ),
    .X(_00761_));
 a22o_1 _19198_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[13] ),
    .A2(net688),
    .B1(net324),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[13] ),
    .X(_00762_));
 mux2_1 _19199_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[14] ),
    .A1(_08393_),
    .S(net711),
    .X(_00763_));
 a22o_1 _19200_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[15] ),
    .A2(net688),
    .B1(net324),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[15] ),
    .X(_00764_));
 mux2_1 _19201_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[16] ),
    .A1(_08311_),
    .S(net713),
    .X(_00765_));
 mux2_1 _19202_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[17] ),
    .A1(_08279_),
    .S(net712),
    .X(_00766_));
 and2_1 _19203_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[18] ),
    .B(net698),
    .X(_04447_));
 a31o_1 _19204_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[2] ),
    .A2(net713),
    .A3(net386),
    .B1(_04447_),
    .X(_00767_));
 a22o_1 _19205_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[19] ),
    .A2(net696),
    .B1(net331),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[3] ),
    .X(_00768_));
 a22o_1 _19206_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[20] ),
    .A2(net698),
    .B1(net333),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[4] ),
    .X(_00769_));
 a22o_1 _19207_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[21] ),
    .A2(net696),
    .B1(net331),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[5] ),
    .X(_00770_));
 a22o_1 _19208_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[22] ),
    .A2(net696),
    .B1(net331),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[6] ),
    .X(_00771_));
 a22o_1 _19209_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[23] ),
    .A2(net690),
    .B1(net327),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ),
    .X(_00772_));
 a22o_1 _19210_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[24] ),
    .A2(net688),
    .B1(net324),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[8] ),
    .X(_00773_));
 a22o_1 _19211_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[25] ),
    .A2(net690),
    .B1(net327),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[9] ),
    .X(_00774_));
 a22o_1 _19212_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[26] ),
    .A2(net688),
    .B1(net325),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[10] ),
    .X(_00775_));
 and2_1 _19213_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[27] ),
    .B(net690),
    .X(_04448_));
 a31o_1 _19214_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[11] ),
    .A2(net710),
    .A3(net373),
    .B1(_04448_),
    .X(_00776_));
 a22o_1 _19215_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[28] ),
    .A2(net690),
    .B1(net327),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[12] ),
    .X(_00777_));
 mux2_1 _19216_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[29] ),
    .A1(_08190_),
    .S(net710),
    .X(_00778_));
 a22o_1 _19217_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[30] ),
    .A2(net690),
    .B1(net327),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[14] ),
    .X(_00779_));
 a22o_1 _19218_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[31] ),
    .A2(net692),
    .B1(net324),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[15] ),
    .X(_00780_));
 a22o_1 _19219_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[32] ),
    .A2(net697),
    .B1(net332),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[0] ),
    .X(_00781_));
 a22o_1 _19220_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[33] ),
    .A2(net694),
    .B1(net332),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[1] ),
    .X(_00782_));
 a22o_1 _19221_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[34] ),
    .A2(net698),
    .B1(net333),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[2] ),
    .X(_00783_));
 a22o_1 _19222_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[35] ),
    .A2(net695),
    .B1(net329),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[3] ),
    .X(_00784_));
 a22o_1 _19223_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[36] ),
    .A2(net693),
    .B1(net329),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[4] ),
    .X(_00785_));
 a22o_1 _19224_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[37] ),
    .A2(net697),
    .B1(net332),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[5] ),
    .X(_00786_));
 mux2_1 _19225_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[38] ),
    .A1(_08208_),
    .S(net712),
    .X(_00787_));
 a22o_1 _19226_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[39] ),
    .A2(net691),
    .B1(net327),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[7] ),
    .X(_00788_));
 a22o_1 _19227_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[40] ),
    .A2(net688),
    .B1(net325),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[8] ),
    .X(_00789_));
 a22o_1 _19228_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[41] ),
    .A2(net690),
    .B1(net328),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[9] ),
    .X(_00790_));
 a22o_1 _19229_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[42] ),
    .A2(net688),
    .B1(net324),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[10] ),
    .X(_00791_));
 a22o_1 _19230_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[43] ),
    .A2(net690),
    .B1(net328),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[11] ),
    .X(_00792_));
 and2_1 _19231_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[44] ),
    .B(net688),
    .X(_04449_));
 a31o_1 _19232_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[12] ),
    .A2(net710),
    .A3(net373),
    .B1(_04449_),
    .X(_00793_));
 a22o_1 _19233_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[45] ),
    .A2(net689),
    .B1(net326),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[13] ),
    .X(_00794_));
 mux2_1 _19234_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[46] ),
    .A1(_08388_),
    .S(net711),
    .X(_00795_));
 a22o_1 _19235_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[47] ),
    .A2(net684),
    .B1(net325),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[15] ),
    .X(_00796_));
 a22o_1 _19236_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[48] ),
    .A2(net697),
    .B1(net332),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[0] ),
    .X(_00797_));
 a22o_1 _19237_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[49] ),
    .A2(net695),
    .B1(net330),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[1] ),
    .X(_00798_));
 a22o_1 _19238_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[50] ),
    .A2(net698),
    .B1(net333),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[2] ),
    .X(_00799_));
 a22o_1 _19239_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[51] ),
    .A2(net693),
    .B1(net330),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[3] ),
    .X(_00800_));
 a22o_1 _19240_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[52] ),
    .A2(net695),
    .B1(net329),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[4] ),
    .X(_00801_));
 a22o_1 _19241_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[53] ),
    .A2(net696),
    .B1(net331),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[5] ),
    .X(_00802_));
 a22o_1 _19242_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[54] ),
    .A2(net693),
    .B1(net329),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[6] ),
    .X(_00803_));
 a22o_1 _19243_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[55] ),
    .A2(net689),
    .B1(net326),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[7] ),
    .X(_00804_));
 a22o_1 _19244_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[56] ),
    .A2(net687),
    .B1(net323),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[8] ),
    .X(_00805_));
 a22o_1 _19245_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[57] ),
    .A2(net689),
    .B1(net326),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[9] ),
    .X(_00806_));
 a22o_1 _19246_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[58] ),
    .A2(net686),
    .B1(net323),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[10] ),
    .X(_00807_));
 a22o_1 _19247_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[59] ),
    .A2(net686),
    .B1(net323),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[11] ),
    .X(_00808_));
 a22o_1 _19248_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[60] ),
    .A2(net686),
    .B1(net323),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[12] ),
    .X(_00809_));
 a22o_1 _19249_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[61] ),
    .A2(net689),
    .B1(net326),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[13] ),
    .X(_00810_));
 a22o_1 _19250_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[62] ),
    .A2(net689),
    .B1(net326),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[14] ),
    .X(_00811_));
 a22o_1 _19251_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[63] ),
    .A2(net685),
    .B1(net322),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[15] ),
    .X(_00812_));
 a22o_1 _19252_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[64] ),
    .A2(net697),
    .B1(net332),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ),
    .X(_00813_));
 and2_1 _19253_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[65] ),
    .B(net694),
    .X(_04450_));
 a31o_1 _19254_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[1] ),
    .A2(net712),
    .A3(net384),
    .B1(_04450_),
    .X(_00814_));
 mux2_1 _19255_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[66] ),
    .A1(_08246_),
    .S(net713),
    .X(_00815_));
 and2_1 _19256_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[67] ),
    .B(net694),
    .X(_04451_));
 a31o_1 _19257_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[3] ),
    .A2(net712),
    .A3(net384),
    .B1(_04451_),
    .X(_00816_));
 mux2_1 _19258_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[68] ),
    .A1(_08160_),
    .S(net713),
    .X(_00817_));
 mux2_1 _19259_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[69] ),
    .A1(_08359_),
    .S(net712),
    .X(_00818_));
 and2_1 _19260_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[70] ),
    .B(net693),
    .X(_04452_));
 a31o_1 _19261_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[6] ),
    .A2(net712),
    .A3(net384),
    .B1(_04452_),
    .X(_00819_));
 a22o_1 _19262_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[71] ),
    .A2(net691),
    .B1(net327),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ),
    .X(_00820_));
 and2_1 _19263_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[72] ),
    .B(net686),
    .X(_04453_));
 a31o_1 _19264_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[8] ),
    .A2(net710),
    .A3(net373),
    .B1(_04453_),
    .X(_00821_));
 and2_1 _19265_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[73] ),
    .B(net689),
    .X(_04454_));
 a31o_1 _19266_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[9] ),
    .A2(net711),
    .A3(net371),
    .B1(_04454_),
    .X(_00822_));
 a22o_1 _19267_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[74] ),
    .A2(net687),
    .B1(net323),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ),
    .X(_00823_));
 and2_1 _19268_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[75] ),
    .B(net686),
    .X(_04455_));
 a31o_1 _19269_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[11] ),
    .A2(net710),
    .A3(net373),
    .B1(_04455_),
    .X(_00824_));
 and2_1 _19270_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[76] ),
    .B(net685),
    .X(_04456_));
 a31o_1 _19271_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[12] ),
    .A2(net710),
    .A3(net373),
    .B1(_04456_),
    .X(_00825_));
 and2_1 _19272_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[77] ),
    .B(net684),
    .X(_04457_));
 a31o_1 _19273_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[13] ),
    .A2(net710),
    .A3(net374),
    .B1(_04457_),
    .X(_00826_));
 and2_1 _19274_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[78] ),
    .B(net684),
    .X(_04458_));
 a31o_1 _19275_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[14] ),
    .A2(net710),
    .A3(net373),
    .B1(_04458_),
    .X(_00827_));
 and2_1 _19276_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[79] ),
    .B(net685),
    .X(_04459_));
 a31o_1 _19277_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[15] ),
    .A2(net710),
    .A3(net374),
    .B1(_04459_),
    .X(_00828_));
 and2_1 _19278_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[80] ),
    .B(net697),
    .X(_04460_));
 a31o_1 _19279_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[0] ),
    .A2(net713),
    .A3(net387),
    .B1(_04460_),
    .X(_00829_));
 a22o_1 _19280_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[81] ),
    .A2(net694),
    .B1(net330),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[1] ),
    .X(_00830_));
 a22o_1 _19281_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[82] ),
    .A2(net698),
    .B1(net333),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[2] ),
    .X(_00831_));
 a22o_1 _19282_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[83] ),
    .A2(net694),
    .B1(net330),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[3] ),
    .X(_00832_));
 a22o_1 _19283_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[84] ),
    .A2(net693),
    .B1(net329),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[4] ),
    .X(_00833_));
 a22o_1 _19284_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[85] ),
    .A2(net695),
    .B1(net330),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[5] ),
    .X(_00834_));
 a22o_1 _19285_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[86] ),
    .A2(net693),
    .B1(net329),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[6] ),
    .X(_00835_));
 a22o_1 _19286_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[87] ),
    .A2(net691),
    .B1(net327),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ),
    .X(_00836_));
 a22o_1 _19287_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[88] ),
    .A2(net686),
    .B1(net323),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[8] ),
    .X(_00837_));
 a22o_1 _19288_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[89] ),
    .A2(net689),
    .B1(net326),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[9] ),
    .X(_00838_));
 and2_1 _19289_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[90] ),
    .B(net687),
    .X(_04461_));
 a31o_1 _19290_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[10] ),
    .A2(net710),
    .A3(net373),
    .B1(_04461_),
    .X(_00839_));
 a22o_1 _19291_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[91] ),
    .A2(net686),
    .B1(net323),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[11] ),
    .X(_00840_));
 a22o_1 _19292_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[92] ),
    .A2(net685),
    .B1(net322),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[12] ),
    .X(_00841_));
 a22o_1 _19293_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[93] ),
    .A2(net684),
    .B1(net322),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[13] ),
    .X(_00842_));
 a22o_1 _19294_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[94] ),
    .A2(net684),
    .B1(net325),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[14] ),
    .X(_00843_));
 a22o_1 _19295_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[95] ),
    .A2(net684),
    .B1(net322),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[15] ),
    .X(_00844_));
 a22o_1 _19296_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[96] ),
    .A2(net696),
    .B1(net331),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[0] ),
    .X(_00845_));
 a22o_1 _19297_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[97] ),
    .A2(net694),
    .B1(net330),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[1] ),
    .X(_00846_));
 a22o_1 _19298_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[98] ),
    .A2(net698),
    .B1(net333),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[2] ),
    .X(_00847_));
 a22o_1 _19299_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[99] ),
    .A2(net694),
    .B1(net330),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[3] ),
    .X(_00848_));
 a22o_1 _19300_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[100] ),
    .A2(net693),
    .B1(net329),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[4] ),
    .X(_00849_));
 and2_1 _19301_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[101] ),
    .B(net694),
    .X(_04462_));
 a31o_1 _19302_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[5] ),
    .A2(net712),
    .A3(net384),
    .B1(_04462_),
    .X(_00850_));
 a22o_1 _19303_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[102] ),
    .A2(net693),
    .B1(net329),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[6] ),
    .X(_00851_));
 a22o_1 _19304_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[103] ),
    .A2(net691),
    .B1(net326),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[7] ),
    .X(_00852_));
 a22o_1 _19305_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[104] ),
    .A2(net686),
    .B1(net323),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[8] ),
    .X(_00853_));
 mux2_1 _19306_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[105] ),
    .A1(_08173_),
    .S(net711),
    .X(_00854_));
 a22o_1 _19307_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[106] ),
    .A2(net687),
    .B1(net324),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ),
    .X(_00855_));
 a22o_1 _19308_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[107] ),
    .A2(net686),
    .B1(net323),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[11] ),
    .X(_00856_));
 a22o_1 _19309_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[108] ),
    .A2(net685),
    .B1(net322),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[12] ),
    .X(_00857_));
 a22o_1 _19310_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[109] ),
    .A2(net689),
    .B1(net326),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[13] ),
    .X(_00858_));
 a22o_1 _19311_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[110] ),
    .A2(net684),
    .B1(net325),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[14] ),
    .X(_00859_));
 a22o_1 _19312_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[111] ),
    .A2(net684),
    .B1(net322),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[15] ),
    .X(_00860_));
 a22o_1 _19313_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[112] ),
    .A2(net697),
    .B1(net332),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[0] ),
    .X(_00861_));
 a22o_1 _19314_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[113] ),
    .A2(net694),
    .B1(net330),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[1] ),
    .X(_00862_));
 a22o_1 _19315_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[114] ),
    .A2(net698),
    .B1(net333),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[2] ),
    .X(_00863_));
 a22o_1 _19316_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[115] ),
    .A2(net694),
    .B1(net330),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[3] ),
    .X(_00864_));
 a22o_1 _19317_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[116] ),
    .A2(net693),
    .B1(net329),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[4] ),
    .X(_00865_));
 and2_1 _19318_ (.A(\digitop_pav2.sec_inst.r128.reg128_o[117] ),
    .B(net695),
    .X(_04463_));
 a31o_1 _19319_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[5] ),
    .A2(net712),
    .A3(net384),
    .B1(_04463_),
    .X(_00866_));
 a22o_1 _19320_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[118] ),
    .A2(net693),
    .B1(net329),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[6] ),
    .X(_00867_));
 a22o_1 _19321_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[119] ),
    .A2(net689),
    .B1(net326),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[7] ),
    .X(_00868_));
 a22o_1 _19322_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[120] ),
    .A2(net686),
    .B1(net323),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[8] ),
    .X(_00869_));
 mux2_1 _19323_ (.A0(\digitop_pav2.sec_inst.r128.reg128_o[121] ),
    .A1(_08172_),
    .S(net711),
    .X(_00870_));
 a22o_1 _19324_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[122] ),
    .A2(net687),
    .B1(net324),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[10] ),
    .X(_00871_));
 a22o_1 _19325_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[123] ),
    .A2(net685),
    .B1(net322),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[11] ),
    .X(_00872_));
 a22o_1 _19326_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[124] ),
    .A2(net685),
    .B1(net322),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[12] ),
    .X(_00873_));
 a22o_1 _19327_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[125] ),
    .A2(net689),
    .B1(net326),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[13] ),
    .X(_00874_));
 a22o_1 _19328_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[126] ),
    .A2(net684),
    .B1(net322),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[14] ),
    .X(_00875_));
 a22o_1 _19329_ (.A1(\digitop_pav2.sec_inst.r128.reg128_o[127] ),
    .A2(net684),
    .B1(net322),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[15] ),
    .X(_00876_));
 or2_2 _19330_ (.A(_08500_),
    .B(_08847_),
    .X(_04464_));
 nor2_2 _19331_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[6] ),
    .B(_04464_),
    .Y(_04465_));
 a21o_1 _19332_ (.A1(\digitop_pav2.sec_inst.shift_out.j_ctr[0] ),
    .A2(_04464_),
    .B1(_04465_),
    .X(_00877_));
 a22o_1 _19333_ (.A1(\digitop_pav2.sec_inst.shift_out.j_ctr[1] ),
    .A2(_04464_),
    .B1(_04465_),
    .B2(\digitop_pav2.sec_inst.shift_out.j_ctr[0] ),
    .X(_00878_));
 a22o_1 _19334_ (.A1(\digitop_pav2.sec_inst.shift_out.j_ctr[2] ),
    .A2(_04464_),
    .B1(_04465_),
    .B2(\digitop_pav2.sec_inst.shift_out.j_ctr[1] ),
    .X(_00879_));
 a22o_1 _19335_ (.A1(\digitop_pav2.sec_inst.shift_out.j_ctr[3] ),
    .A2(_04464_),
    .B1(_04465_),
    .B2(\digitop_pav2.sec_inst.shift_out.j_ctr[2] ),
    .X(_00880_));
 a22o_1 _19336_ (.A1(\digitop_pav2.sec_inst.shift_out.j_ctr[4] ),
    .A2(_04464_),
    .B1(_04465_),
    .B2(\digitop_pav2.sec_inst.shift_out.j_ctr[3] ),
    .X(_00881_));
 a22o_1 _19337_ (.A1(\digitop_pav2.sec_inst.shift_out.j_ctr[5] ),
    .A2(_04464_),
    .B1(_04465_),
    .B2(\digitop_pav2.sec_inst.shift_out.j_ctr[4] ),
    .X(_00882_));
 and2_1 _19338_ (.A(\digitop_pav2.sec_inst.shift_out.j_ctr[6] ),
    .B(_04464_),
    .X(_04466_));
 a21o_1 _19339_ (.A1(\digitop_pav2.sec_inst.shift_out.j_ctr[5] ),
    .A2(_04465_),
    .B1(_04466_),
    .X(_00883_));
 mux2_1 _19340_ (.A0(\digitop_pav2.sec_inst.shift_in.s9.q[0] ),
    .A1(net1641),
    .S(net590),
    .X(_00884_));
 mux2_1 _19341_ (.A0(\digitop_pav2.sec_inst.shift_in.s9.q[1] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s9.q[0] ),
    .S(net590),
    .X(_00885_));
 mux2_1 _19342_ (.A0(\digitop_pav2.sec_inst.shift_in.s9.q[2] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s9.q[1] ),
    .S(net590),
    .X(_00886_));
 mux2_1 _19343_ (.A0(\digitop_pav2.sec_inst.shift_in.s9.q[3] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s9.q[2] ),
    .S(net590),
    .X(_00887_));
 mux2_1 _19344_ (.A0(\digitop_pav2.sec_inst.shift_in.s9.q[4] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s9.q[3] ),
    .S(net590),
    .X(_00888_));
 mux2_1 _19345_ (.A0(\digitop_pav2.sec_inst.shift_in.s9.q[5] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s9.q[4] ),
    .S(net590),
    .X(_00889_));
 mux2_1 _19346_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[30] ),
    .A1(\digitop_pav2.sec_inst.shift_in.s9.q[5] ),
    .S(_03018_),
    .X(_00890_));
 mux2_1 _19347_ (.A0(\digitop_pav2.sec_inst.ld_r.reg96_i[31] ),
    .A1(\digitop_pav2.sec_inst.ld_r.reg96_i[30] ),
    .S(net590),
    .X(_00891_));
 or4b_1 _19348_ (.A(\digitop_pav2.sec_inst.shift_out.st[4] ),
    .B(\digitop_pav2.sec_inst.shift_out.st[7] ),
    .C(\digitop_pav2.sec_inst.shift_out.st[0] ),
    .D_N(\digitop_pav2.sec_inst.shift_out.ctr[0] ),
    .X(_04467_));
 xnor2_1 _19349_ (.A(\digitop_pav2.sec_inst.shift_out.ctr[0] ),
    .B(_08493_),
    .Y(_00892_));
 xnor2_1 _19350_ (.A(\digitop_pav2.sec_inst.shift_out.ctr[1] ),
    .B(_04467_),
    .Y(_00893_));
 nor2_1 _19351_ (.A(_08493_),
    .B(_08498_),
    .Y(_04468_));
 o21ba_1 _19352_ (.A1(_08493_),
    .A2(_08497_),
    .B1_N(net706),
    .X(_04469_));
 nor2_1 _19353_ (.A(_04468_),
    .B(_04469_),
    .Y(_00894_));
 mux2_1 _19354_ (.A0(net704),
    .A1(_08495_),
    .S(_04468_),
    .X(_00895_));
 a21o_1 _19355_ (.A1(net712),
    .A2(net1653),
    .B1(net702),
    .X(_00896_));
 and2_1 _19356_ (.A(_10855_),
    .B(_10857_),
    .X(_00897_));
 and3_1 _19357_ (.A(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[1] ),
    .B(_01284_),
    .C(_10857_),
    .X(_00898_));
 nor2_1 _19358_ (.A(_07063_),
    .B(_03662_),
    .Y(_04470_));
 nor2_1 _19359_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[9] ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.state[2] ),
    .Y(_04471_));
 or4_1 _19360_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.state[9] ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.state[2] ),
    .C(\digitop_pav2.invent_inst.invent_sel_pav2.state[7] ),
    .D(\digitop_pav2.invent_inst.invent_sel_pav2.state[11] ),
    .X(_04472_));
 o22a_1 _19361_ (.A1(_07909_),
    .A2(_10330_),
    .B1(_04472_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.state[1] ),
    .X(_04473_));
 o31a_1 _19362_ (.A1(_07892_),
    .A2(_07900_),
    .A3(_04471_),
    .B1(_04470_),
    .X(_04474_));
 and4bb_1 _19363_ (.A_N(\digitop_pav2.access_inst.access_ctrl0.nvm_busy_i ),
    .B_N(_10562_),
    .C(_04473_),
    .D(_04474_),
    .X(_04475_));
 mux2_1 _19364_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[0] ),
    .A1(net1135),
    .S(net158),
    .X(_00899_));
 mux2_1 _19365_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[1] ),
    .A1(net1133),
    .S(net158),
    .X(_00900_));
 mux2_1 _19366_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[2] ),
    .A1(net1129),
    .S(net157),
    .X(_00901_));
 mux2_1 _19367_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[3] ),
    .A1(net1125),
    .S(net157),
    .X(_00902_));
 mux2_1 _19368_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[4] ),
    .A1(net1122),
    .S(net157),
    .X(_00903_));
 mux2_1 _19369_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[5] ),
    .A1(net1119),
    .S(net157),
    .X(_00904_));
 mux2_1 _19370_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[6] ),
    .A1(net1116),
    .S(net158),
    .X(_00905_));
 mux2_1 _19371_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[7] ),
    .A1(net1113),
    .S(net157),
    .X(_00906_));
 mux2_1 _19372_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[8] ),
    .A1(net1109),
    .S(net157),
    .X(_00907_));
 mux2_1 _19373_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[9] ),
    .A1(net1105),
    .S(net158),
    .X(_00908_));
 mux2_1 _19374_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[10] ),
    .A1(net1101),
    .S(net158),
    .X(_00909_));
 mux2_1 _19375_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[11] ),
    .A1(net1097),
    .S(net157),
    .X(_00910_));
 mux2_1 _19376_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[12] ),
    .A1(net1095),
    .S(net158),
    .X(_00911_));
 mux2_1 _19377_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[13] ),
    .A1(net1092),
    .S(net157),
    .X(_00912_));
 mux2_1 _19378_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[14] ),
    .A1(net1088),
    .S(net157),
    .X(_00913_));
 mux2_1 _19379_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[15] ),
    .A1(net1085),
    .S(net157),
    .X(_00914_));
 and2_1 _19380_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.timeout_en_t1 ),
    .B(_10315_),
    .X(_04476_));
 xor2_1 _19381_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[0] ),
    .B(_04476_),
    .X(_00915_));
 and4_1 _19382_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[0] ),
    .B(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[1] ),
    .C(\digitop_pav2.proc_ctrl_inst.cmdfsm.timeout_en_t1 ),
    .D(_10315_),
    .X(_04477_));
 a21oi_1 _19383_ (.A1(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[0] ),
    .A2(_04476_),
    .B1(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[1] ),
    .Y(_04478_));
 nor2_1 _19384_ (.A(_04477_),
    .B(_04478_),
    .Y(_00916_));
 xor2_1 _19385_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[2] ),
    .B(_04477_),
    .X(_00917_));
 and3_1 _19386_ (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[2] ),
    .B(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[3] ),
    .C(_04477_),
    .X(_04479_));
 a21o_1 _19387_ (.A1(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[2] ),
    .A2(_04477_),
    .B1(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[3] ),
    .X(_04480_));
 and2b_1 _19388_ (.A_N(_04479_),
    .B(_04480_),
    .X(_00918_));
 xnor2_1 _19389_ (.A(_07158_),
    .B(_04479_),
    .Y(_00919_));
 xnor2_1 _19390_ (.A(\digitop_pav2.func_rng_data[5] ),
    .B(\digitop_pav2.func_rng_data[8] ),
    .Y(_04481_));
 xnor2_1 _19391_ (.A(\digitop_pav2.func_rng_data[7] ),
    .B(\digitop_pav2.func_rng_data[9] ),
    .Y(_04482_));
 nor2_1 _19392_ (.A(_04481_),
    .B(_04482_),
    .Y(_04483_));
 a211o_1 _19393_ (.A1(_04481_),
    .A2(_04482_),
    .B1(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[0] ),
    .C1(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[1] ),
    .X(_04484_));
 xnor2_1 _19394_ (.A(\digitop_pav2.func_rng_data[3] ),
    .B(\digitop_pav2.func_rng_data[8] ),
    .Y(_04485_));
 xnor2_1 _19395_ (.A(\digitop_pav2.func_rng_data[5] ),
    .B(\digitop_pav2.func_rng_data[11] ),
    .Y(_04486_));
 xnor2_1 _19396_ (.A(_04485_),
    .B(_04486_),
    .Y(_04487_));
 or4bb_1 _19397_ (.A(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[1] ),
    .B(_04487_),
    .C_N(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[0] ),
    .D_N(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[2] ),
    .X(_04488_));
 nand2b_1 _19398_ (.A_N(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[2] ),
    .B(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[0] ),
    .Y(_04489_));
 or2_1 _19399_ (.A(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[1] ),
    .B(_04489_),
    .X(_04490_));
 nand2_1 _19400_ (.A(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[1] ),
    .B(_04489_),
    .Y(_04491_));
 nand2_1 _19401_ (.A(_04490_),
    .B(_04491_),
    .Y(_04492_));
 o211a_1 _19402_ (.A1(_04481_),
    .A2(_04489_),
    .B1(_04490_),
    .C1(_04491_),
    .X(_04493_));
 or4b_1 _19403_ (.A(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[0] ),
    .B(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[1] ),
    .C(_04485_),
    .D_N(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[2] ),
    .X(_04494_));
 o311a_1 _19404_ (.A1(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[2] ),
    .A2(_04483_),
    .A3(_04484_),
    .B1(_04493_),
    .C1(_04494_),
    .X(_04495_));
 xnor2_1 _19405_ (.A(\digitop_pav2.func_rng_data[8] ),
    .B(\digitop_pav2.func_rng_data[9] ),
    .Y(_04496_));
 mux2_1 _19406_ (.A0(_04496_),
    .A1(_04485_),
    .S(_04490_),
    .X(_04497_));
 and2_1 _19407_ (.A(\digitop_pav2.func_rng_data[11] ),
    .B(_04497_),
    .X(_04498_));
 o21ai_1 _19408_ (.A1(\digitop_pav2.func_rng_data[11] ),
    .A2(_04497_),
    .B1(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[0] ),
    .Y(_04499_));
 xnor2_1 _19409_ (.A(\digitop_pav2.func_rng_data[7] ),
    .B(\digitop_pav2.func_rng_data[8] ),
    .Y(_04500_));
 and3b_1 _19410_ (.A_N(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[0] ),
    .B(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[2] ),
    .C(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[1] ),
    .X(_04501_));
 mux2_1 _19411_ (.A0(\digitop_pav2.func_rng_data[9] ),
    .A1(\digitop_pav2.func_rng_data[11] ),
    .S(_04501_),
    .X(_04502_));
 xnor2_1 _19412_ (.A(_04500_),
    .B(_04502_),
    .Y(_04503_));
 o22a_1 _19413_ (.A1(_04498_),
    .A2(_04499_),
    .B1(_04503_),
    .B2(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[0] ),
    .X(_04504_));
 xnor2_1 _19414_ (.A(\digitop_pav2.func_rng_data[13] ),
    .B(_04504_),
    .Y(_04505_));
 a22o_1 _19415_ (.A1(_04488_),
    .A2(_04495_),
    .B1(_04505_),
    .B2(_04492_),
    .X(_04506_));
 nor2_1 _19416_ (.A(\digitop_pav2.func_rng_data[14] ),
    .B(\digitop_pav2.func_rng_data[15] ),
    .Y(_04507_));
 or4_1 _19417_ (.A(\digitop_pav2.func_rng_data[10] ),
    .B(\digitop_pav2.func_rng_data[11] ),
    .C(\digitop_pav2.func_rng_data[12] ),
    .D(\digitop_pav2.func_rng_data[13] ),
    .X(_04508_));
 or4_1 _19418_ (.A(\digitop_pav2.func_rng_data[3] ),
    .B(\digitop_pav2.func_rng_data[4] ),
    .C(\digitop_pav2.func_rng_data[6] ),
    .D(\digitop_pav2.func_rng_data[7] ),
    .X(_04509_));
 or4_1 _19419_ (.A(\digitop_pav2.func_rng_data[5] ),
    .B(\digitop_pav2.func_rng_data[0] ),
    .C(\digitop_pav2.func_rng_data[1] ),
    .D(\digitop_pav2.func_rng_data[2] ),
    .X(_04510_));
 or3_1 _19420_ (.A(\digitop_pav2.func_rng_data[8] ),
    .B(\digitop_pav2.func_rng_data[9] ),
    .C(_04510_),
    .X(_04511_));
 o31a_1 _19421_ (.A1(_04508_),
    .A2(_04509_),
    .A3(_04511_),
    .B1(_04507_),
    .X(_04512_));
 a21oi_1 _19422_ (.A1(\digitop_pav2.func_rng_data[14] ),
    .A2(\digitop_pav2.func_rng_data[15] ),
    .B1(_04512_),
    .Y(_04513_));
 xnor2_1 _19423_ (.A(_04506_),
    .B(_04513_),
    .Y(_04514_));
 mux2_1 _19424_ (.A0(\digitop_pav2.func_rng_data[0] ),
    .A1(_04514_),
    .S(net678),
    .X(_00920_));
 mux2_1 _19425_ (.A0(\digitop_pav2.func_rng_data[1] ),
    .A1(\digitop_pav2.func_rng_data[0] ),
    .S(net678),
    .X(_00921_));
 mux2_1 _19426_ (.A0(\digitop_pav2.func_rng_data[2] ),
    .A1(\digitop_pav2.func_rng_data[1] ),
    .S(net679),
    .X(_00922_));
 mux2_1 _19427_ (.A0(\digitop_pav2.func_rng_data[3] ),
    .A1(\digitop_pav2.func_rng_data[2] ),
    .S(net678),
    .X(_00923_));
 mux2_1 _19428_ (.A0(\digitop_pav2.func_rng_data[4] ),
    .A1(\digitop_pav2.func_rng_data[3] ),
    .S(net679),
    .X(_00924_));
 mux2_1 _19429_ (.A0(\digitop_pav2.func_rng_data[5] ),
    .A1(\digitop_pav2.func_rng_data[4] ),
    .S(net679),
    .X(_00925_));
 mux2_1 _19430_ (.A0(\digitop_pav2.func_rng_data[6] ),
    .A1(\digitop_pav2.func_rng_data[5] ),
    .S(net678),
    .X(_00926_));
 mux2_1 _19431_ (.A0(\digitop_pav2.func_rng_data[7] ),
    .A1(\digitop_pav2.func_rng_data[6] ),
    .S(net678),
    .X(_00927_));
 mux2_1 _19432_ (.A0(\digitop_pav2.func_rng_data[8] ),
    .A1(\digitop_pav2.func_rng_data[7] ),
    .S(net679),
    .X(_00928_));
 mux2_1 _19433_ (.A0(\digitop_pav2.func_rng_data[9] ),
    .A1(\digitop_pav2.func_rng_data[8] ),
    .S(net679),
    .X(_00929_));
 mux2_1 _19434_ (.A0(\digitop_pav2.func_rng_data[10] ),
    .A1(\digitop_pav2.func_rng_data[9] ),
    .S(net678),
    .X(_00930_));
 mux2_1 _19435_ (.A0(\digitop_pav2.func_rng_data[11] ),
    .A1(\digitop_pav2.func_rng_data[10] ),
    .S(net678),
    .X(_00931_));
 mux2_1 _19436_ (.A0(\digitop_pav2.func_rng_data[12] ),
    .A1(\digitop_pav2.func_rng_data[11] ),
    .S(net678),
    .X(_00932_));
 mux2_1 _19437_ (.A0(\digitop_pav2.func_rng_data[13] ),
    .A1(\digitop_pav2.func_rng_data[12] ),
    .S(net679),
    .X(_00933_));
 mux2_1 _19438_ (.A0(\digitop_pav2.func_rng_data[14] ),
    .A1(\digitop_pav2.func_rng_data[13] ),
    .S(net678),
    .X(_00934_));
 mux2_1 _19439_ (.A0(\digitop_pav2.func_rng_data[15] ),
    .A1(\digitop_pav2.func_rng_data[14] ),
    .S(net678),
    .X(_00935_));
 nand2_1 _19440_ (.A(_07316_),
    .B(_09146_),
    .Y(_04515_));
 a21oi_1 _19441_ (.A1(_10484_),
    .A2(_04515_),
    .B1(_10315_),
    .Y(_04516_));
 and3_1 _19442_ (.A(_07330_),
    .B(net1229),
    .C(_10498_),
    .X(_04517_));
 a31o_1 _19443_ (.A1(net1292),
    .A2(_07276_),
    .A3(net1162),
    .B1(_10481_),
    .X(_04518_));
 o21ai_1 _19444_ (.A1(_07312_),
    .A2(_07352_),
    .B1(_07299_),
    .Y(_04519_));
 a21o_1 _19445_ (.A1(net1181),
    .A2(_07347_),
    .B1(_08518_),
    .X(_04520_));
 or2_1 _19446_ (.A(_07354_),
    .B(_04520_),
    .X(_04521_));
 o21a_1 _19447_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[12] ),
    .A2(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[3] ),
    .B1(net156),
    .X(_04522_));
 a221o_1 _19448_ (.A1(_07283_),
    .A2(_09034_),
    .B1(_10459_),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[5] ),
    .C1(_04522_),
    .X(_04523_));
 or2_1 _19449_ (.A(_09013_),
    .B(_10496_),
    .X(_04524_));
 or4_1 _19450_ (.A(_07327_),
    .B(_07348_),
    .C(_09019_),
    .D(_09024_),
    .X(_04525_));
 or4_1 _19451_ (.A(net1295),
    .B(_10505_),
    .C(_04524_),
    .D(_04525_),
    .X(_04526_));
 or4_1 _19452_ (.A(_04519_),
    .B(_04521_),
    .C(_04523_),
    .D(_04526_),
    .X(_04527_));
 or4_1 _19453_ (.A(_10876_),
    .B(_04517_),
    .C(_04518_),
    .D(_04527_),
    .X(_04528_));
 or3b_1 _19454_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[1] ),
    .B(net1287),
    .C_N(_04528_),
    .X(_04529_));
 nand2_1 _19455_ (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[1] ),
    .B(_10315_),
    .Y(_04530_));
 o311a_1 _19456_ (.A1(_07087_),
    .A2(_09032_),
    .A3(_04516_),
    .B1(_04529_),
    .C1(_04530_),
    .X(_04531_));
 a21o_1 _19457_ (.A1(net1286),
    .A2(_04516_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[1] ),
    .X(_04532_));
 mux2_1 _19458_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.en_i ),
    .A1(_04532_),
    .S(_04531_),
    .X(_00936_));
 nor2_1 _19459_ (.A(_07242_),
    .B(net1219),
    .Y(_04533_));
 or2_1 _19460_ (.A(_07066_),
    .B(_07303_),
    .X(_04534_));
 a31o_1 _19461_ (.A1(_07242_),
    .A2(_07307_),
    .A3(_04534_),
    .B1(_07245_),
    .X(_04535_));
 or3_1 _19462_ (.A(net1253),
    .B(net1219),
    .C(_07263_),
    .X(_04536_));
 o21a_1 _19463_ (.A1(net1232),
    .A2(_07286_),
    .B1(_04536_),
    .X(_04537_));
 or2_1 _19464_ (.A(net1232),
    .B(_07263_),
    .X(_04538_));
 nor2_1 _19465_ (.A(_07249_),
    .B(_04538_),
    .Y(_04539_));
 or3_1 _19466_ (.A(net1232),
    .B(_07241_),
    .C(net1230),
    .X(_04540_));
 o21ai_1 _19467_ (.A1(net1219),
    .A2(_07280_),
    .B1(_04540_),
    .Y(_04541_));
 nor2_1 _19468_ (.A(_04539_),
    .B(_04541_),
    .Y(_04542_));
 inv_2 _19469_ (.A(_04542_),
    .Y(_04543_));
 nor2_1 _19470_ (.A(_07242_),
    .B(net1231),
    .Y(_04544_));
 or4_1 _19471_ (.A(_07247_),
    .B(net1196),
    .C(_09030_),
    .D(_04544_),
    .X(_04545_));
 nand2_1 _19472_ (.A(net1232),
    .B(net1231),
    .Y(_04546_));
 a22o_1 _19473_ (.A1(_07065_),
    .A2(_07268_),
    .B1(_04546_),
    .B2(_07251_),
    .X(_04547_));
 nor2_1 _19474_ (.A(_07239_),
    .B(_07255_),
    .Y(_04548_));
 nor2_1 _19475_ (.A(net1232),
    .B(_07303_),
    .Y(_04549_));
 and3b_1 _19476_ (.A_N(_07263_),
    .B(_07065_),
    .C(_07249_),
    .X(_04550_));
 or3_1 _19477_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[5] ),
    .B(_07250_),
    .C(_07263_),
    .X(_04551_));
 or4_1 _19478_ (.A(net1186),
    .B(_04548_),
    .C(_04549_),
    .D(_04550_),
    .X(_04552_));
 or4_1 _19479_ (.A(_07295_),
    .B(_07331_),
    .C(_04547_),
    .D(_04552_),
    .X(_04553_));
 nor2_1 _19480_ (.A(_04545_),
    .B(_04553_),
    .Y(_04554_));
 and4_1 _19481_ (.A(_04535_),
    .B(_04537_),
    .C(_04542_),
    .D(_04554_),
    .X(_04555_));
 nor2_1 _19482_ (.A(_04539_),
    .B(_04547_),
    .Y(_04556_));
 a21oi_1 _19483_ (.A1(_04535_),
    .A2(_04556_),
    .B1(_07071_),
    .Y(_04557_));
 a21o_1 _19484_ (.A1(_07071_),
    .A2(_04544_),
    .B1(_07292_),
    .X(_04558_));
 or4_1 _19485_ (.A(net1196),
    .B(_04541_),
    .C(_04555_),
    .D(_04558_),
    .X(_04559_));
 a311o_1 _19486_ (.A1(net1252),
    .A2(_07899_),
    .A3(_04550_),
    .B1(_04557_),
    .C1(_04559_),
    .X(_04560_));
 nand2_1 _19487_ (.A(net1322),
    .B(net1030),
    .Y(_04561_));
 nor3_1 _19488_ (.A(_07262_),
    .B(_07263_),
    .C(net1230),
    .Y(_04562_));
 a31o_1 _19489_ (.A1(net1297),
    .A2(_04561_),
    .A3(_04562_),
    .B1(net1197),
    .X(_04563_));
 a41o_1 _19490_ (.A1(\digitop_pav2.proc_ctrl_inst.cmd.state[5] ),
    .A2(net1252),
    .A3(_07071_),
    .A4(_07308_),
    .B1(_04563_),
    .X(_04564_));
 a31o_1 _19491_ (.A1(net1298),
    .A2(_07287_),
    .A3(_07308_),
    .B1(_04564_),
    .X(_04565_));
 or4_1 _19492_ (.A(_07067_),
    .B(net1231),
    .C(_07286_),
    .D(_04561_),
    .X(_04566_));
 o21ai_1 _19493_ (.A1(net1297),
    .A2(_04566_),
    .B1(_07265_),
    .Y(_04567_));
 a21oi_1 _19494_ (.A1(_07066_),
    .A2(_04549_),
    .B1(_04544_),
    .Y(_04568_));
 a21o_1 _19495_ (.A1(_07309_),
    .A2(_04534_),
    .B1(net1219),
    .X(_04569_));
 o31a_1 _19496_ (.A1(net1254),
    .A2(net1231),
    .A3(_07286_),
    .B1(_04569_),
    .X(_04570_));
 or3_1 _19497_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[1] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state[0] ),
    .C(_04538_),
    .X(_04571_));
 nor3b_1 _19498_ (.A(_07246_),
    .B(net1231),
    .C_N(net1230),
    .Y(_04572_));
 nor2_1 _19499_ (.A(_04533_),
    .B(_04572_),
    .Y(_04573_));
 o2111a_1 _19500_ (.A1(net1219),
    .A2(_07286_),
    .B1(_04571_),
    .C1(_04573_),
    .D1(_07071_),
    .X(_04574_));
 a22o_1 _19501_ (.A1(net1297),
    .A2(_04568_),
    .B1(_04570_),
    .B2(_04574_),
    .X(_04575_));
 and3_1 _19502_ (.A(net1252),
    .B(net1030),
    .C(_04550_),
    .X(_04576_));
 or3_1 _19503_ (.A(_07241_),
    .B(net1231),
    .C(net1230),
    .X(_04577_));
 o22a_1 _19504_ (.A1(_07241_),
    .A2(_07266_),
    .B1(_07303_),
    .B2(_07065_),
    .X(_04578_));
 or3b_1 _19505_ (.A(net1297),
    .B(_04578_),
    .C_N(net1252),
    .X(_04579_));
 nand2_1 _19506_ (.A(_04577_),
    .B(_04579_),
    .Y(_04580_));
 or3b_1 _19507_ (.A(net1198),
    .B(net1187),
    .C_N(_04536_),
    .X(_04581_));
 or3_1 _19508_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[5] ),
    .B(net1298),
    .C(_07267_),
    .X(_04582_));
 nand2_1 _19509_ (.A(_07257_),
    .B(_04582_),
    .Y(_04583_));
 or4_1 _19510_ (.A(net1185),
    .B(_04580_),
    .C(_04581_),
    .D(_04583_),
    .X(_04584_));
 or4b_1 _19511_ (.A(_04567_),
    .B(_04584_),
    .C(_04576_),
    .D_N(_04575_),
    .X(_04585_));
 nor2_1 _19512_ (.A(_04565_),
    .B(_04585_),
    .Y(_04586_));
 inv_2 _19513_ (.A(_04586_),
    .Y(_04587_));
 and2_2 _19514_ (.A(net1304),
    .B(_10461_),
    .X(_04588_));
 nand2b_1 _19515_ (.A_N(_04560_),
    .B(_04588_),
    .Y(_04589_));
 nor2_1 _19516_ (.A(_04586_),
    .B(_04589_),
    .Y(_04590_));
 nor2_1 _19517_ (.A(_07067_),
    .B(_04537_),
    .Y(_04591_));
 or3_1 _19518_ (.A(_07240_),
    .B(_07246_),
    .C(_07262_),
    .X(_04592_));
 or3_1 _19519_ (.A(_07067_),
    .B(_07241_),
    .C(_07288_),
    .X(_04593_));
 o211a_1 _19520_ (.A1(_04534_),
    .A2(_04546_),
    .B1(_04592_),
    .C1(_04593_),
    .X(_04594_));
 or3b_1 _19521_ (.A(net1297),
    .B(_04533_),
    .C_N(_04594_),
    .X(_04595_));
 o21a_1 _19522_ (.A1(net1254),
    .A2(_04537_),
    .B1(_04577_),
    .X(_04596_));
 o2bb2a_1 _19523_ (.A1_N(net1297),
    .A2_N(_04596_),
    .B1(_04595_),
    .B2(_04591_),
    .X(_04597_));
 or4_1 _19524_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[5] ),
    .B(net1298),
    .C(_07241_),
    .D(net1230),
    .X(_04598_));
 and4_1 _19525_ (.A(net1297),
    .B(_07249_),
    .C(_07253_),
    .D(_07287_),
    .X(_04599_));
 a31o_1 _19526_ (.A1(net1253),
    .A2(net1297),
    .A3(_04549_),
    .B1(_04599_),
    .X(_04600_));
 or3b_1 _19527_ (.A(_07292_),
    .B(_04600_),
    .C_N(_04598_),
    .X(_04601_));
 or4_1 _19528_ (.A(net1298),
    .B(net1232),
    .C(_07246_),
    .D(_07250_),
    .X(_04602_));
 o21ai_1 _19529_ (.A1(\digitop_pav2.proc_ctrl_inst.cmd.state[4] ),
    .A2(_04551_),
    .B1(_04602_),
    .Y(_04603_));
 or4_1 _19530_ (.A(net1195),
    .B(_04548_),
    .C(_04601_),
    .D(_04603_),
    .X(_04604_));
 or4_1 _19531_ (.A(net1187),
    .B(_04576_),
    .C(_04583_),
    .D(_04604_),
    .X(_04605_));
 or3_2 _19532_ (.A(_04565_),
    .B(_04597_),
    .C(_04605_),
    .X(_04606_));
 a2111o_1 _19533_ (.A1(net1322),
    .A2(_07067_),
    .B1(_07241_),
    .C1(_07288_),
    .D1(\digitop_pav2.proc_ctrl_inst.cmd.state[1] ),
    .X(_04607_));
 o221a_1 _19534_ (.A1(net1231),
    .A2(_07280_),
    .B1(_04538_),
    .B2(_07066_),
    .C1(_04607_),
    .X(_04608_));
 a31o_1 _19535_ (.A1(_04570_),
    .A2(_04596_),
    .A3(_04608_),
    .B1(net1297),
    .X(_04609_));
 nand2_1 _19536_ (.A(_04582_),
    .B(_04602_),
    .Y(_04610_));
 or4_1 _19537_ (.A(net1186),
    .B(net1195),
    .C(_04591_),
    .D(_04610_),
    .X(_04611_));
 or4b_1 _19538_ (.A(_04545_),
    .B(_04601_),
    .C(_04611_),
    .D_N(_04609_),
    .X(_04612_));
 or2_1 _19539_ (.A(_04565_),
    .B(_04612_),
    .X(_04613_));
 inv_2 _19540_ (.A(_04613_),
    .Y(_04614_));
 nor2_1 _19541_ (.A(_04606_),
    .B(_04614_),
    .Y(_04615_));
 a21o_1 _19542_ (.A1(_07071_),
    .A2(_04576_),
    .B1(_07252_),
    .X(_04616_));
 o21ai_1 _19543_ (.A1(\digitop_pav2.proc_ctrl_inst.cmd.state[5] ),
    .A2(_07267_),
    .B1(_07304_),
    .Y(_04617_));
 a211o_1 _19544_ (.A1(_04546_),
    .A2(_04617_),
    .B1(_04572_),
    .C1(_04543_),
    .X(_04618_));
 mux2_1 _19545_ (.A0(_04548_),
    .A1(_04618_),
    .S(_07071_),
    .X(_04619_));
 or4_1 _19546_ (.A(_07361_),
    .B(_04581_),
    .C(_04603_),
    .D(_04619_),
    .X(_04620_));
 or4_2 _19547_ (.A(_04564_),
    .B(_04567_),
    .C(_04616_),
    .D(_04620_),
    .X(_04621_));
 inv_2 _19548_ (.A(_04621_),
    .Y(_04622_));
 o21bai_1 _19549_ (.A1(\digitop_pav2.proc_ctrl_inst.cmd.state[4] ),
    .A2(_04551_),
    .B1_N(_04591_),
    .Y(_04623_));
 or2_1 _19550_ (.A(_07280_),
    .B(_07288_),
    .X(_04624_));
 and4bb_1 _19551_ (.A_N(_04541_),
    .B_N(_04548_),
    .C(_04593_),
    .D(_04624_),
    .X(_04625_));
 a21oi_1 _19552_ (.A1(_04573_),
    .A2(_04625_),
    .B1(net1298),
    .Y(_04626_));
 or3_1 _19553_ (.A(_04544_),
    .B(_04549_),
    .C(_04610_),
    .X(_04627_));
 or4_1 _19554_ (.A(_07260_),
    .B(net1185),
    .C(_07361_),
    .D(_04580_),
    .X(_04628_));
 a211o_1 _19555_ (.A1(net1297),
    .A2(_04623_),
    .B1(_04626_),
    .C1(_04628_),
    .X(_04629_));
 or3_1 _19556_ (.A(_04563_),
    .B(_04627_),
    .C(_04629_),
    .X(_04630_));
 nor2_1 _19557_ (.A(_04616_),
    .B(_04630_),
    .Y(_04631_));
 nor2_1 _19558_ (.A(_04622_),
    .B(_04631_),
    .Y(_04632_));
 a21o_1 _19559_ (.A1(net1241),
    .A2(_10695_),
    .B1(_09096_),
    .X(_04633_));
 a41o_1 _19560_ (.A1(_04590_),
    .A2(_04615_),
    .A3(_04632_),
    .A4(_04633_),
    .B1(net1281),
    .X(_00937_));
 nor2_1 _19561_ (.A(_04587_),
    .B(_04589_),
    .Y(_04634_));
 nor2_1 _19562_ (.A(_04621_),
    .B(_04630_),
    .Y(_04635_));
 and2_1 _19563_ (.A(_04606_),
    .B(_04613_),
    .X(_04636_));
 a41o_1 _19564_ (.A1(_10911_),
    .A2(_04634_),
    .A3(_04635_),
    .A4(_04636_),
    .B1(net1280),
    .X(_00938_));
 nor2_1 _19565_ (.A(_04621_),
    .B(_04631_),
    .Y(_04637_));
 nor2_1 _19566_ (.A(_04606_),
    .B(_04613_),
    .Y(_04638_));
 a41o_1 _19567_ (.A1(_10911_),
    .A2(_04590_),
    .A3(_04637_),
    .A4(_04638_),
    .B1(net1277),
    .X(_00939_));
 and3_1 _19568_ (.A(_04590_),
    .B(_04606_),
    .C(_04614_),
    .X(_04639_));
 a41o_1 _19569_ (.A1(net1241),
    .A2(_09096_),
    .A3(_04635_),
    .A4(_04639_),
    .B1(\digitop_pav2.access_inst.access_check0.g_write_i ),
    .X(_00940_));
 a31o_1 _19570_ (.A1(_04632_),
    .A2(_04634_),
    .A3(_04638_),
    .B1(net1275),
    .X(_00941_));
 and3_1 _19571_ (.A(_04560_),
    .B(_04586_),
    .C(_04588_),
    .X(_04640_));
 a31o_1 _19572_ (.A1(_04632_),
    .A2(_04636_),
    .A3(_04640_),
    .B1(net1273),
    .X(_00942_));
 a41o_1 _19573_ (.A1(_10903_),
    .A2(_04615_),
    .A3(_04634_),
    .A4(_04637_),
    .B1(net1267),
    .X(_00943_));
 o21a_1 _19574_ (.A1(\digitop_pav2.pie_inst.fsm.past_ctr[4] ),
    .A2(_09578_),
    .B1(net495),
    .X(_04641_));
 o2111a_1 _19575_ (.A1(net493),
    .A2(_04641_),
    .B1(_09649_),
    .C1(_09581_),
    .D1(_09585_),
    .X(_00944_));
 a41o_1 _19576_ (.A1(_10912_),
    .A2(_04615_),
    .A3(_04635_),
    .A4(_04640_),
    .B1(\digitop_pav2.access_inst.access_check0.g_propwrite_i ),
    .X(_00945_));
 a31o_1 _19577_ (.A1(_09096_),
    .A2(_04632_),
    .A3(_04639_),
    .B1(net1263),
    .X(_00946_));
 nand2_1 _19578_ (.A(_04588_),
    .B(_04631_),
    .Y(_04642_));
 nor2_1 _19579_ (.A(_04622_),
    .B(_04642_),
    .Y(_04643_));
 a41o_1 _19580_ (.A1(_09096_),
    .A2(_04560_),
    .A3(_04638_),
    .A4(_04643_),
    .B1(net1258),
    .X(_00947_));
 and4_1 _19581_ (.A(_10883_),
    .B(_04560_),
    .C(_04587_),
    .D(_04588_),
    .X(_04644_));
 a31o_1 _19582_ (.A1(_04632_),
    .A2(_04636_),
    .A3(_04644_),
    .B1(\digitop_pav2.proc_ctrl_inst.cmd.g_sec_auth_o ),
    .X(_00948_));
 or4_1 _19583_ (.A(\digitop_pav2.proc_ctrl_inst.ebv.state[8] ),
    .B(\digitop_pav2.proc_ctrl_inst.ebv.state[1] ),
    .C(\digitop_pav2.proc_ctrl_inst.ebv.state[3] ),
    .D(\digitop_pav2.proc_ctrl_inst.ebv.state[7] ),
    .X(_04645_));
 or4_1 _19584_ (.A(\digitop_pav2.proc_ctrl_inst.ebv.state[6] ),
    .B(\digitop_pav2.proc_ctrl_inst.ebv.state[11] ),
    .C(\digitop_pav2.proc_ctrl_inst.ebv.state[13] ),
    .D(_04645_),
    .X(_04646_));
 a31o_1 _19585_ (.A1(net1299),
    .A2(net970),
    .A3(_04646_),
    .B1(\digitop_pav2.proc_ctrl_inst.ebv.invalid ),
    .X(_00949_));
 a31o_1 _19586_ (.A1(\digitop_pav2.proc_ctrl_inst.profsm.r1_ff ),
    .A2(_07161_),
    .A3(net969),
    .B1(_10902_),
    .X(_04647_));
 nor2_1 _19587_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[2] ),
    .B(_04647_),
    .Y(_04648_));
 a22o_1 _19588_ (.A1(\digitop_pav2.proc_ctrl_inst.profsm.r1_rise_ff ),
    .A2(_10902_),
    .B1(_04648_),
    .B2(_10878_),
    .X(_00955_));
 mux2_1 _19589_ (.A0(net1254),
    .A1(_04613_),
    .S(_04588_),
    .X(_00957_));
 mux2_1 _19590_ (.A0(net1253),
    .A1(_04606_),
    .S(_04588_),
    .X(_00958_));
 o21a_1 _19591_ (.A1(\digitop_pav2.proc_ctrl_inst.cmd.state[2] ),
    .A2(_04588_),
    .B1(_04642_),
    .X(_00959_));
 mux2_1 _19592_ (.A0(\digitop_pav2.proc_ctrl_inst.cmd.state[3] ),
    .A1(_04621_),
    .S(_04588_),
    .X(_00960_));
 mux2_1 _19593_ (.A0(net1252),
    .A1(_04587_),
    .S(_04588_),
    .X(_00961_));
 o21a_1 _19594_ (.A1(\digitop_pav2.proc_ctrl_inst.cmd.state[5] ),
    .A2(_04588_),
    .B1(_04589_),
    .X(_00962_));
 nor2_1 _19595_ (.A(net1396),
    .B(net968),
    .Y(_00224_));
 nand2_1 _19596_ (.A(net1245),
    .B(_10879_),
    .Y(_04649_));
 a41o_1 _19597_ (.A1(net1246),
    .A2(_09031_),
    .A3(net1163),
    .A4(_10879_),
    .B1(_10884_),
    .X(_04650_));
 a21oi_1 _19598_ (.A1(_08871_),
    .A2(_10883_),
    .B1(net1196),
    .Y(_04651_));
 or3_1 _19599_ (.A(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[1] ),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[0] ),
    .C(_07161_),
    .X(_04652_));
 a211oi_2 _19600_ (.A1(_08870_),
    .A2(_09143_),
    .B1(_04651_),
    .C1(_04652_),
    .Y(_04653_));
 or3_1 _19601_ (.A(_10908_),
    .B(_10911_),
    .C(_04649_),
    .X(_04654_));
 o2111ai_4 _19602_ (.A1(_10906_),
    .A2(_10911_),
    .B1(_04650_),
    .C1(_04653_),
    .D1(_04654_),
    .Y(_04655_));
 nor2_2 _19603_ (.A(_10884_),
    .B(net528),
    .Y(_04656_));
 or2_2 _19604_ (.A(_10884_),
    .B(net528),
    .X(_04657_));
 nand2_1 _19605_ (.A(_08877_),
    .B(_04656_),
    .Y(_04658_));
 a21bo_1 _19606_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[0] ),
    .A2(net527),
    .B1_N(_04658_),
    .X(_00975_));
 nand2_1 _19607_ (.A(_08889_),
    .B(_04656_),
    .Y(_04659_));
 a21bo_1 _19608_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[1] ),
    .A2(net527),
    .B1_N(_04659_),
    .X(_00976_));
 nand2_1 _19609_ (.A(_08891_),
    .B(_04656_),
    .Y(_04660_));
 a21bo_1 _19610_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[2] ),
    .A2(net528),
    .B1_N(_04660_),
    .X(_00977_));
 nand2_1 _19611_ (.A(\digitop_pav2.access_inst.access_transceiver0.handle_i[3] ),
    .B(net528),
    .Y(_04661_));
 o21ai_1 _19612_ (.A1(_08887_),
    .A2(_04657_),
    .B1(_04661_),
    .Y(_00978_));
 nand2_1 _19613_ (.A(_08890_),
    .B(_04656_),
    .Y(_04662_));
 a21bo_1 _19614_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[4] ),
    .A2(net528),
    .B1_N(_04662_),
    .X(_00979_));
 nand2_1 _19615_ (.A(\digitop_pav2.access_inst.access_transceiver0.handle_i[5] ),
    .B(net527),
    .Y(_04663_));
 o21ai_1 _19616_ (.A1(_08896_),
    .A2(_04657_),
    .B1(_04663_),
    .Y(_00980_));
 nand2_1 _19617_ (.A(\digitop_pav2.access_inst.access_transceiver0.handle_i[6] ),
    .B(net527),
    .Y(_04664_));
 o21ai_1 _19618_ (.A1(_08901_),
    .A2(_04657_),
    .B1(_04664_),
    .Y(_00981_));
 nand2_1 _19619_ (.A(\digitop_pav2.access_inst.access_transceiver0.handle_i[7] ),
    .B(net527),
    .Y(_04665_));
 o21ai_1 _19620_ (.A1(_08898_),
    .A2(_04657_),
    .B1(_04665_),
    .Y(_00982_));
 nand2_1 _19621_ (.A(\digitop_pav2.access_inst.access_transceiver0.handle_i[8] ),
    .B(net528),
    .Y(_04666_));
 o21ai_1 _19622_ (.A1(_08904_),
    .A2(_04657_),
    .B1(_04666_),
    .Y(_00983_));
 nor2_1 _19623_ (.A(_08912_),
    .B(_04657_),
    .Y(_04667_));
 a21o_1 _19624_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[9] ),
    .A2(net527),
    .B1(_04667_),
    .X(_00984_));
 nand2_1 _19625_ (.A(_08908_),
    .B(_04656_),
    .Y(_04668_));
 a21bo_1 _19626_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[10] ),
    .A2(net528),
    .B1_N(_04668_),
    .X(_00985_));
 nand2_1 _19627_ (.A(_08913_),
    .B(_04656_),
    .Y(_04669_));
 a21bo_1 _19628_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[11] ),
    .A2(net527),
    .B1_N(_04669_),
    .X(_00986_));
 nand2_1 _19629_ (.A(_08909_),
    .B(_04656_),
    .Y(_04670_));
 a21bo_1 _19630_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[12] ),
    .A2(net528),
    .B1_N(_04670_),
    .X(_00987_));
 nand2_1 _19631_ (.A(\digitop_pav2.access_inst.access_transceiver0.handle_i[13] ),
    .B(net527),
    .Y(_04671_));
 a21bo_1 _19632_ (.A1(_08883_),
    .A2(_04656_),
    .B1_N(_04671_),
    .X(_00988_));
 nand2_1 _19633_ (.A(_08881_),
    .B(_04656_),
    .Y(_04672_));
 a21bo_1 _19634_ (.A1(\digitop_pav2.access_inst.access_transceiver0.handle_i[14] ),
    .A2(net527),
    .B1_N(_04672_),
    .X(_00989_));
 nand2_1 _19635_ (.A(\digitop_pav2.access_inst.access_transceiver0.handle_i[15] ),
    .B(net527),
    .Y(_04673_));
 o21ai_1 _19636_ (.A1(_08879_),
    .A2(_04657_),
    .B1(_04673_),
    .Y(_00990_));
 nand2b_1 _19637_ (.A_N(_10981_),
    .B(_11002_),
    .Y(_04674_));
 nor2_1 _19638_ (.A(\digitop_pav2.pie_inst.fsm.state[1] ),
    .B(_10990_),
    .Y(_04675_));
 o32ai_4 _19639_ (.A1(\digitop_pav2.pie_inst.fsm.state[1] ),
    .A2(_10990_),
    .A3(_04674_),
    .B1(_10981_),
    .B2(\digitop_pav2.pie_inst.fsm.state[0] ),
    .Y(_00991_));
 nand2_1 _19640_ (.A(\digitop_pav2.pie_inst.fsm.state[0] ),
    .B(_04675_),
    .Y(_04676_));
 a32o_1 _19641_ (.A1(\digitop_pav2.pie_inst.fsm.state[0] ),
    .A2(_04674_),
    .A3(_04675_),
    .B1(_10991_),
    .B2(_10992_),
    .X(_00992_));
 nor2_1 _19642_ (.A(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[4] ),
    .B(_08874_),
    .Y(_04677_));
 xor2_1 _19643_ (.A(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[2] ),
    .B(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[3] ),
    .X(_04678_));
 xnor2_1 _19644_ (.A(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[1] ),
    .B(_04678_),
    .Y(_04679_));
 a22o_1 _19645_ (.A1(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[0] ),
    .A2(_08874_),
    .B1(_04677_),
    .B2(_04679_),
    .X(_00993_));
 a21oi_1 _19646_ (.A1(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[0] ),
    .A2(_04678_),
    .B1(_08512_),
    .Y(_04680_));
 a22o_1 _19647_ (.A1(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[1] ),
    .A2(_08874_),
    .B1(_04677_),
    .B2(_04680_),
    .X(_00994_));
 mux2_1 _19648_ (.A0(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[2] ),
    .A1(_07118_),
    .S(_08882_),
    .X(_04681_));
 a22o_1 _19649_ (.A1(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[2] ),
    .A2(_08874_),
    .B1(_04677_),
    .B2(_04681_),
    .X(_00995_));
 a31o_1 _19650_ (.A1(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[2] ),
    .A2(_08512_),
    .A3(_08873_),
    .B1(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[3] ),
    .X(_04682_));
 o31a_1 _19651_ (.A1(_07119_),
    .A2(_08514_),
    .A3(_08874_),
    .B1(_04682_),
    .X(_00996_));
 mux2_1 _19652_ (.A0(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[4] ),
    .A1(_08514_),
    .S(_08873_),
    .X(_00997_));
 o31a_1 _19653_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[7] ),
    .A2(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[6] ),
    .A3(net1293),
    .B1(net1250),
    .X(_04683_));
 o211a_1 _19654_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.timeout_en_t1 ),
    .A2(_04683_),
    .B1(_07070_),
    .C1(_07150_),
    .X(_00999_));
 or3b_1 _19655_ (.A(_09140_),
    .B(_04520_),
    .C_N(_10545_),
    .X(_04684_));
 or3_1 _19656_ (.A(_07354_),
    .B(_04517_),
    .C(_04524_),
    .X(_04685_));
 or3b_1 _19657_ (.A(_10485_),
    .B(_04522_),
    .C_N(_10543_),
    .X(_04686_));
 or3_1 _19658_ (.A(_07317_),
    .B(_04525_),
    .C(_04686_),
    .X(_04687_));
 a21o_1 _19659_ (.A1(net1288),
    .A2(net1186),
    .B1(_10505_),
    .X(_04688_));
 a211o_1 _19660_ (.A1(_07313_),
    .A2(_07351_),
    .B1(_04687_),
    .C1(_04688_),
    .X(_04689_));
 or4_1 _19661_ (.A(_09011_),
    .B(_04684_),
    .C(_04685_),
    .D(_04689_),
    .X(_04690_));
 or2_1 _19662_ (.A(_10873_),
    .B(_04518_),
    .X(_04691_));
 or3_1 _19663_ (.A(_10500_),
    .B(_10874_),
    .C(_04518_),
    .X(_04692_));
 or3_1 _19664_ (.A(_10511_),
    .B(_04690_),
    .C(_04692_),
    .X(_04693_));
 nor2_1 _19665_ (.A(_08488_),
    .B(_10519_),
    .Y(_04694_));
 a221o_1 _19666_ (.A1(_09153_),
    .A2(_10523_),
    .B1(_04694_),
    .B2(_07278_),
    .C1(_04693_),
    .X(_04695_));
 a211o_1 _19667_ (.A1(_07325_),
    .A2(_09029_),
    .B1(net1187),
    .C1(_07070_),
    .X(_04696_));
 a2bb2o_1 _19668_ (.A1_N(_04693_),
    .A2_N(_04696_),
    .B1(_04695_),
    .B2(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmd_abort_b ),
    .X(_01000_));
 nand2_1 _19669_ (.A(\digitop_pav2.proc_ctrl_inst.inst_checker.state[9] ),
    .B(net1167),
    .Y(_04697_));
 a31o_1 _19670_ (.A1(net1304),
    .A2(_07275_),
    .A3(_04697_),
    .B1(_10519_),
    .X(_04698_));
 a21oi_1 _19671_ (.A1(_07257_),
    .A2(_07265_),
    .B1(_07279_),
    .Y(_04699_));
 or4_1 _19672_ (.A(_09019_),
    .B(_10499_),
    .C(_04517_),
    .D(_04699_),
    .X(_04700_));
 a32o_1 _19673_ (.A1(net1305),
    .A2(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[7] ),
    .A3(net1195),
    .B1(_07363_),
    .B2(net1218),
    .X(_04701_));
 a21o_1 _19674_ (.A1(net1288),
    .A2(_07302_),
    .B1(_10531_),
    .X(_04702_));
 or4_1 _19675_ (.A(_07327_),
    .B(_07348_),
    .C(_09024_),
    .D(_04522_),
    .X(_04703_));
 or4_1 _19676_ (.A(_07354_),
    .B(_09141_),
    .C(_10505_),
    .D(_04702_),
    .X(_04704_));
 or4_1 _19677_ (.A(_07328_),
    .B(_09013_),
    .C(_10496_),
    .D(_04703_),
    .X(_04705_));
 or4_1 _19678_ (.A(_10522_),
    .B(_10532_),
    .C(_04701_),
    .D(_04705_),
    .X(_04706_));
 or3_1 _19679_ (.A(_10452_),
    .B(_04704_),
    .C(_04706_),
    .X(_04707_));
 a211o_1 _19680_ (.A1(_07292_),
    .A2(_07363_),
    .B1(_07365_),
    .C1(_07318_),
    .X(_04708_));
 a31o_1 _19681_ (.A1(net1294),
    .A2(_07259_),
    .A3(net1183),
    .B1(_04708_),
    .X(_04709_));
 and3_1 _19682_ (.A(net1292),
    .B(_07269_),
    .C(_07276_),
    .X(_04710_));
 a2111o_1 _19683_ (.A1(net1198),
    .A2(_07278_),
    .B1(_10524_),
    .C1(_04684_),
    .D1(_04707_),
    .X(_04711_));
 a2111o_1 _19684_ (.A1(net1291),
    .A2(_10527_),
    .B1(_04700_),
    .C1(_04709_),
    .D1(_04710_),
    .X(_04712_));
 or3_1 _19685_ (.A(_04691_),
    .B(_04711_),
    .C(_04712_),
    .X(_04713_));
 a311o_1 _19686_ (.A1(net1293),
    .A2(net1186),
    .A3(_04698_),
    .B1(_04713_),
    .C1(_09128_),
    .X(_04714_));
 nand2_1 _19687_ (.A(_07299_),
    .B(_09017_),
    .Y(_04715_));
 a31o_1 _19688_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[1] ),
    .A2(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[0] ),
    .A3(_09015_),
    .B1(net1250),
    .X(_04716_));
 a22o_1 _19689_ (.A1(net1295),
    .A2(_07310_),
    .B1(_04715_),
    .B2(_04716_),
    .X(_04717_));
 or3_1 _19690_ (.A(_07363_),
    .B(_10510_),
    .C(_04717_),
    .X(_04718_));
 mux2_1 _19691_ (.A0(_04718_),
    .A1(net1250),
    .S(_04714_),
    .X(_01001_));
 o221a_1 _19692_ (.A1(_07258_),
    .A2(_07260_),
    .B1(_07325_),
    .B2(_07259_),
    .C1(net1294),
    .X(_04719_));
 or3_1 _19693_ (.A(\digitop_pav2.pie_inst.delend_o ),
    .B(_07366_),
    .C(_04688_),
    .X(_04720_));
 or4_1 _19694_ (.A(_10513_),
    .B(_04687_),
    .C(_04719_),
    .D(_04720_),
    .X(_04721_));
 or4b_1 _19695_ (.A(_04520_),
    .B(_04685_),
    .C(_04721_),
    .D_N(_10545_),
    .X(_04722_));
 nor2_1 _19696_ (.A(_04692_),
    .B(_04722_),
    .Y(_04723_));
 o221a_1 _19697_ (.A1(_07259_),
    .A2(_07270_),
    .B1(_10519_),
    .B2(net1249),
    .C1(_07278_),
    .X(_04724_));
 o32a_1 _19698_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdctr.cmdctr_end3 ),
    .A2(net1249),
    .A3(net1189),
    .B1(_07298_),
    .B2(_07284_),
    .X(_04725_));
 o21a_1 _19699_ (.A1(net1249),
    .A2(_09152_),
    .B1(_10523_),
    .X(_04726_));
 a21o_1 _19700_ (.A1(net1305),
    .A2(net1187),
    .B1(net1195),
    .X(_04727_));
 o311a_1 _19701_ (.A1(net1249),
    .A2(_07306_),
    .A3(net1189),
    .B1(net1229),
    .C1(_07313_),
    .X(_04728_));
 a311o_1 _19702_ (.A1(net1295),
    .A2(net1184),
    .A3(_04727_),
    .B1(_04728_),
    .C1(_07328_),
    .X(_04729_));
 or4_1 _19703_ (.A(_10452_),
    .B(_04725_),
    .C(_04726_),
    .D(_04729_),
    .X(_04730_));
 a211o_1 _19704_ (.A1(_07278_),
    .A2(_10869_),
    .B1(_04724_),
    .C1(_04730_),
    .X(_04731_));
 mux2_1 _19705_ (.A0(net1249),
    .A1(_04731_),
    .S(_04723_),
    .X(_01002_));
 or2_1 _19706_ (.A(_04521_),
    .B(_04710_),
    .X(_04732_));
 nor2_1 _19707_ (.A(_04699_),
    .B(_04732_),
    .Y(_04733_));
 inv_2 _19708_ (.A(_04733_),
    .Y(_04734_));
 and2b_1 _19709_ (.A_N(_09131_),
    .B(_07284_),
    .X(_04735_));
 or4b_1 _19710_ (.A(_09018_),
    .B(_04702_),
    .C(_04735_),
    .D_N(_10545_),
    .X(_04736_));
 or4_1 _19711_ (.A(_04517_),
    .B(_04526_),
    .C(_04686_),
    .D(_04736_),
    .X(_04737_));
 a21o_1 _19712_ (.A1(_07298_),
    .A2(_09138_),
    .B1(_04737_),
    .X(_04738_));
 a21oi_1 _19713_ (.A1(net1291),
    .A2(_10527_),
    .B1(_04738_),
    .Y(_04739_));
 o211a_1 _19714_ (.A1(_07248_),
    .A2(_07279_),
    .B1(_04733_),
    .C1(_04739_),
    .X(_04740_));
 nor4b_1 _19715_ (.A(_10499_),
    .B(_10512_),
    .C(_04691_),
    .D_N(_04740_),
    .Y(_04741_));
 a311o_1 _19716_ (.A1(net1245),
    .A2(_09153_),
    .A3(_10523_),
    .B1(_04519_),
    .C1(_10510_),
    .X(_04742_));
 mux2_1 _19717_ (.A0(net1244),
    .A1(_04742_),
    .S(_04741_),
    .X(_01003_));
 a21oi_4 _19718_ (.A1(_08870_),
    .A2(_09149_),
    .B1(_07329_),
    .Y(_04743_));
 mux2_1 _19719_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[0] ),
    .A1(\digitop_pav2.memctrl_inst.extra_dt_i[12] ),
    .S(net1022),
    .X(_01004_));
 mux2_1 _19720_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[1] ),
    .A1(\digitop_pav2.memctrl_inst.extra_dt_i[13] ),
    .S(net1022),
    .X(_01005_));
 mux2_1 _19721_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[2] ),
    .A1(\digitop_pav2.memctrl_inst.extra_dt_i[14] ),
    .S(net1022),
    .X(_01006_));
 mux2_1 _19722_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[3] ),
    .A1(\digitop_pav2.memctrl_inst.extra_dt_i[15] ),
    .S(_04743_),
    .X(_01007_));
 mux2_1 _19723_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[4] ),
    .A1(\digitop_pav2.pie_inst.fsm.trcal[4] ),
    .S(net1022),
    .X(_01008_));
 mux2_1 _19724_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[5] ),
    .A1(\digitop_pav2.pie_inst.fsm.trcal[5] ),
    .S(net1022),
    .X(_01009_));
 mux2_1 _19725_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[6] ),
    .A1(\digitop_pav2.pie_inst.fsm.trcal[6] ),
    .S(net1022),
    .X(_01010_));
 mux2_1 _19726_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[7] ),
    .A1(\digitop_pav2.pie_inst.fsm.trcal[7] ),
    .S(_04743_),
    .X(_01011_));
 mux2_1 _19727_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[8] ),
    .A1(\digitop_pav2.pie_inst.fsm.trcal[8] ),
    .S(_04743_),
    .X(_01012_));
 mux2_1 _19728_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[9] ),
    .A1(\digitop_pav2.pie_inst.fsm.trcal[9] ),
    .S(_04743_),
    .X(_01013_));
 mux2_1 _19729_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_trext ),
    .A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[3] ),
    .S(net1022),
    .X(_01014_));
 mux2_1 _19730_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_m[0] ),
    .A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[2] ),
    .S(net1022),
    .X(_01015_));
 mux2_1 _19731_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_m[1] ),
    .A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[1] ),
    .S(net1022),
    .X(_01016_));
 mux2_1 _19732_ (.A0(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_dr ),
    .A1(\digitop_pav2.dr ),
    .S(net1022),
    .X(_01017_));
 nand2_1 _19733_ (.A(_07153_),
    .B(_10449_),
    .Y(_04744_));
 mux2_1 _19734_ (.A0(net1299),
    .A1(\digitop_pav2.fg_tc ),
    .S(_04744_),
    .X(_01018_));
 or4_1 _19735_ (.A(_07284_),
    .B(_07318_),
    .C(_07328_),
    .D(_10496_),
    .X(_04745_));
 a211o_1 _19736_ (.A1(_07260_),
    .A2(_07278_),
    .B1(_04688_),
    .C1(_04745_),
    .X(_04746_));
 a21oi_1 _19737_ (.A1(net1216),
    .A2(_07311_),
    .B1(_07352_),
    .Y(_04747_));
 or2_1 _19738_ (.A(_07298_),
    .B(_04747_),
    .X(_04748_));
 nand2_1 _19739_ (.A(_09017_),
    .B(_10545_),
    .Y(_04749_));
 or2_1 _19740_ (.A(_09013_),
    .B(_04749_),
    .X(_04750_));
 or4_1 _19741_ (.A(net1291),
    .B(net1289),
    .C(net1292),
    .D(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[5] ),
    .X(_04751_));
 or3_1 _19742_ (.A(net1290),
    .B(_10533_),
    .C(_04751_),
    .X(_04752_));
 nor2_1 _19743_ (.A(net1294),
    .B(_04752_),
    .Y(_04753_));
 or4_1 _19744_ (.A(_07317_),
    .B(_07348_),
    .C(_04750_),
    .D(_04753_),
    .X(_04754_));
 or3_1 _19745_ (.A(_04521_),
    .B(_04748_),
    .C(_04754_),
    .X(_04755_));
 or3_2 _19746_ (.A(_04699_),
    .B(_04746_),
    .C(_04755_),
    .X(_04756_));
 nor2_1 _19747_ (.A(_10490_),
    .B(_04756_),
    .Y(_04757_));
 o211a_1 _19748_ (.A1(net1289),
    .A2(_07278_),
    .B1(net1197),
    .C1(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_cgen.fg_tc_rx_i ),
    .X(_04758_));
 or2_1 _19749_ (.A(_09024_),
    .B(_04756_),
    .X(_04759_));
 o22a_1 _19750_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_cgen.fg_tc_rx_i ),
    .A2(_04757_),
    .B1(_04758_),
    .B2(_04759_),
    .X(_01019_));
 nor2_1 _19751_ (.A(_10449_),
    .B(_04756_),
    .Y(_04760_));
 o211a_1 _19752_ (.A1(net1289),
    .A2(_07278_),
    .B1(net1197),
    .C1(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_cgen.en_g_sec_i ),
    .X(_04761_));
 o22a_1 _19753_ (.A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_cgen.en_g_sec_i ),
    .A2(_04760_),
    .B1(_04761_),
    .B2(_04759_),
    .X(_01020_));
 or4_1 _19754_ (.A(_07317_),
    .B(_09024_),
    .C(_10508_),
    .D(_10522_),
    .X(_04762_));
 a2111o_1 _19755_ (.A1(_07310_),
    .A2(_07363_),
    .B1(_04701_),
    .C1(_04753_),
    .D1(_04762_),
    .X(_04763_));
 or4_1 _19756_ (.A(_07298_),
    .B(_04746_),
    .C(_04750_),
    .D(_04763_),
    .X(_04764_));
 nor4_1 _19757_ (.A(_04691_),
    .B(_04700_),
    .C(_04732_),
    .D(_04764_),
    .Y(_04765_));
 and3_1 _19758_ (.A(_07295_),
    .B(_07364_),
    .C(_04765_),
    .X(_04766_));
 o2bb2a_1 _19759_ (.A1_N(_04752_),
    .A2_N(_04765_),
    .B1(_04766_),
    .B2(net973),
    .X(_01021_));
 o31a_1 _19760_ (.A1(_07294_),
    .A2(_07352_),
    .A3(net1189),
    .B1(_04752_),
    .X(_04767_));
 or3b_1 _19761_ (.A(_04749_),
    .B(_04762_),
    .C_N(_04767_),
    .X(_04768_));
 or4_1 _19762_ (.A(_10874_),
    .B(_04746_),
    .C(_04748_),
    .D(_04768_),
    .X(_04769_));
 or4_1 _19763_ (.A(_04517_),
    .B(_04518_),
    .C(_04734_),
    .D(_04769_),
    .X(_04770_));
 nor4_1 _19764_ (.A(_07041_),
    .B(_07294_),
    .C(_10533_),
    .D(_04751_),
    .Y(_04771_));
 mux2_1 _19765_ (.A0(_04771_),
    .A1(\digitop_pav2.proc_ctrl_inst.cmdfsm.ebv_en ),
    .S(_04770_),
    .X(_01022_));
 and4_1 _19766_ (.A(_07130_),
    .B(net969),
    .C(_10892_),
    .D(_10905_),
    .X(_04772_));
 inv_2 _19767_ (.A(_04772_),
    .Y(_04773_));
 and2_1 _19768_ (.A(_09148_),
    .B(_09149_),
    .X(_04774_));
 o2bb2a_1 _19769_ (.A1_N(_07361_),
    .A2_N(_04774_),
    .B1(_09149_),
    .B2(_07312_),
    .X(_04775_));
 o31a_1 _19770_ (.A1(\digitop_pav2.proc_ctrl_inst.profsm.r1_ff ),
    .A2(_09143_),
    .A3(_09151_),
    .B1(_04775_),
    .X(_04776_));
 o221a_1 _19771_ (.A1(\digitop_pav2.proc_ctrl_inst.profsm.r1_ff ),
    .A2(_10484_),
    .B1(_10886_),
    .B2(_04776_),
    .C1(net1246),
    .X(_04777_));
 o21ba_1 _19772_ (.A1(_10887_),
    .A2(_04777_),
    .B1_N(_10882_),
    .X(_04778_));
 o21ai_1 _19773_ (.A1(\digitop_pav2.proc_ctrl_inst.int_pass_t2_flag ),
    .A2(_07305_),
    .B1(_04774_),
    .Y(_04779_));
 or4b_1 _19774_ (.A(net969),
    .B(\digitop_pav2.proc_ctrl_inst.profsm.skip_abort ),
    .C(_09151_),
    .D_N(\digitop_pav2.proc_ctrl_inst.int_pass_t2_flag ),
    .X(_04780_));
 o21a_1 _19775_ (.A1(_07312_),
    .A2(_04779_),
    .B1(_04780_),
    .X(_04781_));
 a21o_1 _19776_ (.A1(net1215),
    .A2(_07312_),
    .B1(_09149_),
    .X(_04782_));
 a311oi_1 _19777_ (.A1(_10879_),
    .A2(_04781_),
    .A3(_04782_),
    .B1(_10896_),
    .C1(net1233),
    .Y(_04783_));
 o31a_1 _19778_ (.A1(\digitop_pav2.proc_ctrl_inst.int_timeout_t2 ),
    .A2(_10894_),
    .A3(_04783_),
    .B1(_10698_),
    .X(_04784_));
 nor2_1 _19779_ (.A(net1215),
    .B(_10879_),
    .Y(_04785_));
 a21o_1 _19780_ (.A1(_07248_),
    .A2(net1215),
    .B1(_10879_),
    .X(_04786_));
 o21a_1 _19781_ (.A1(_10878_),
    .A2(_04775_),
    .B1(_04786_),
    .X(_04787_));
 o311a_1 _19782_ (.A1(net1233),
    .A2(\digitop_pav2.proc_ctrl_inst.int_timeout_t2 ),
    .A3(_04787_),
    .B1(_10695_),
    .C1(net1241),
    .X(_04788_));
 or4_1 _19783_ (.A(_07292_),
    .B(_09149_),
    .C(_10911_),
    .D(_04649_),
    .X(_04789_));
 a311o_1 _19784_ (.A1(net1245),
    .A2(_07361_),
    .A3(_09148_),
    .B1(_10880_),
    .C1(_10904_),
    .X(_04790_));
 o211ai_1 _19785_ (.A1(_09031_),
    .A2(_10877_),
    .B1(_04789_),
    .C1(_04790_),
    .Y(_04791_));
 or3_1 _19786_ (.A(_07248_),
    .B(_07899_),
    .C(_10881_),
    .X(_04792_));
 or3_1 _19787_ (.A(net1215),
    .B(_09149_),
    .C(_04649_),
    .X(_04793_));
 a31o_1 _19788_ (.A1(_10892_),
    .A2(_04792_),
    .A3(_04793_),
    .B1(_10884_),
    .X(_04794_));
 or4b_1 _19789_ (.A(_04772_),
    .B(_04788_),
    .C(_04791_),
    .D_N(_04794_),
    .X(_04795_));
 o32a_1 _19790_ (.A1(_04778_),
    .A2(_04784_),
    .A3(_04795_),
    .B1(_04773_),
    .B2(net1241),
    .X(_01024_));
 o21a_1 _19791_ (.A1(net1216),
    .A2(_09149_),
    .B1(_04775_),
    .X(_04796_));
 nor2_1 _19792_ (.A(_10878_),
    .B(_04796_),
    .Y(_04797_));
 a31o_1 _19793_ (.A1(net1198),
    .A2(_10697_),
    .A3(_10878_),
    .B1(_04797_),
    .X(_04798_));
 o21ai_1 _19794_ (.A1(_04649_),
    .A2(_04781_),
    .B1(_10695_),
    .Y(_04799_));
 a2111o_1 _19795_ (.A1(net1246),
    .A2(_04798_),
    .B1(_04799_),
    .C1(\digitop_pav2.proc_ctrl_inst.int_timeout_t2 ),
    .D1(_10894_),
    .X(_04800_));
 o221a_1 _19796_ (.A1(net1215),
    .A2(_10884_),
    .B1(_10903_),
    .B2(_07289_),
    .C1(_10904_),
    .X(_04801_));
 or3_1 _19797_ (.A(net1233),
    .B(\digitop_pav2.proc_ctrl_inst.profsm.r1_ff ),
    .C(_10484_),
    .X(_04802_));
 o2bb2a_1 _19798_ (.A1_N(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[1] ),
    .A2_N(_04772_),
    .B1(_04801_),
    .B2(_10881_),
    .X(_04803_));
 o211ai_1 _19799_ (.A1(_10882_),
    .A2(_04802_),
    .B1(_04803_),
    .C1(_04800_),
    .Y(_01025_));
 o21ai_1 _19800_ (.A1(_04785_),
    .A2(_04797_),
    .B1(net1246),
    .Y(_04804_));
 or3_1 _19801_ (.A(net1234),
    .B(_10886_),
    .C(_04796_),
    .X(_04805_));
 a32o_1 _19802_ (.A1(_10693_),
    .A2(_04802_),
    .A3(_04805_),
    .B1(_10880_),
    .B2(_09144_),
    .X(_04806_));
 and4_1 _19803_ (.A(net1246),
    .B(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[0] ),
    .C(_07130_),
    .D(_10695_),
    .X(_04807_));
 and3_1 _19804_ (.A(net1198),
    .B(_10878_),
    .C(_04807_),
    .X(_04808_));
 a41o_1 _19805_ (.A1(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[0] ),
    .A2(_09031_),
    .A3(_09096_),
    .A4(_04806_),
    .B1(_04808_),
    .X(_04809_));
 a32o_1 _19806_ (.A1(_10883_),
    .A2(_10892_),
    .A3(_04804_),
    .B1(_04809_),
    .B2(_04773_),
    .X(_04810_));
 a21o_1 _19807_ (.A1(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[2] ),
    .A2(_04772_),
    .B1(_04810_),
    .X(_01026_));
 nand2_1 _19808_ (.A(\digitop_pav2.proc_ctrl_inst.profsm.skip_abort ),
    .B(_04647_),
    .Y(_04811_));
 o21ai_1 _19809_ (.A1(_10463_),
    .A2(_04647_),
    .B1(_04811_),
    .Y(_01027_));
 o2bb2a_1 _19810_ (.A1_N(_07160_),
    .A2_N(_10902_),
    .B1(_04647_),
    .B2(_09146_),
    .X(_01028_));
 nand2_1 _19811_ (.A(\digitop_pav2.pie_inst.fsm.state[1] ),
    .B(_10990_),
    .Y(_04812_));
 a41o_1 _19812_ (.A1(_07145_),
    .A2(\digitop_pav2.pie_inst.delend_o ),
    .A3(_10981_),
    .A4(_04812_),
    .B1(net475),
    .X(_01029_));
 or4_4 _19813_ (.A(net1399),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.piex_dt_rx_done ),
    .C(_11002_),
    .D(_04676_),
    .X(_04813_));
 mux2_1 _19814_ (.A0(\digitop_pav2.pie_inst.fsm.dif_pos_fix[0] ),
    .A1(\digitop_pav2.memctrl_inst.extra_dt_i[12] ),
    .S(_04813_),
    .X(_01030_));
 mux2_1 _19815_ (.A0(\digitop_pav2.pie_inst.fsm.dif_pos_fix[1] ),
    .A1(\digitop_pav2.memctrl_inst.extra_dt_i[13] ),
    .S(_04813_),
    .X(_01031_));
 mux2_1 _19816_ (.A0(\digitop_pav2.pie_inst.fsm.dif_pos_fix[2] ),
    .A1(\digitop_pav2.memctrl_inst.extra_dt_i[14] ),
    .S(_04813_),
    .X(_01032_));
 mux2_1 _19817_ (.A0(\digitop_pav2.pie_inst.fsm.dif_pos_fix[3] ),
    .A1(\digitop_pav2.memctrl_inst.extra_dt_i[15] ),
    .S(_04813_),
    .X(_01033_));
 mux2_1 _19818_ (.A0(\digitop_pav2.pie_inst.fsm.dif_pos_fix[4] ),
    .A1(\digitop_pav2.pie_inst.fsm.trcal[4] ),
    .S(_04813_),
    .X(_01034_));
 mux2_1 _19819_ (.A0(\digitop_pav2.pie_inst.fsm.dif_pos_fix[5] ),
    .A1(\digitop_pav2.pie_inst.fsm.trcal[5] ),
    .S(_04813_),
    .X(_01035_));
 mux2_1 _19820_ (.A0(\digitop_pav2.pie_inst.fsm.dif_pos_fix[6] ),
    .A1(\digitop_pav2.pie_inst.fsm.trcal[6] ),
    .S(_04813_),
    .X(_01036_));
 mux2_1 _19821_ (.A0(\digitop_pav2.pie_inst.fsm.dif_pos_fix[7] ),
    .A1(\digitop_pav2.pie_inst.fsm.trcal[7] ),
    .S(_04813_),
    .X(_01037_));
 mux2_1 _19822_ (.A0(\digitop_pav2.pie_inst.fsm.dif_pos_fix[8] ),
    .A1(\digitop_pav2.pie_inst.fsm.trcal[8] ),
    .S(_04813_),
    .X(_01038_));
 mux2_1 _19823_ (.A0(\digitop_pav2.pie_inst.fsm.dif_pos_fix[9] ),
    .A1(\digitop_pav2.pie_inst.fsm.trcal[9] ),
    .S(_04813_),
    .X(_01039_));
 mux2_1 _19824_ (.A0(\digitop_pav2.memctrl_inst.addr_to_reram[0] ),
    .A1(net1764),
    .S(_07931_),
    .X(_01040_));
 nor2_1 _19825_ (.A(net1753),
    .B(_07925_),
    .Y(_04814_));
 mux2_1 _19826_ (.A0(\digitop_pav2.memctrl_inst.addr_to_reram[1] ),
    .A1(net1754),
    .S(_07931_),
    .X(_01041_));
 o21a_1 _19827_ (.A1(_07922_),
    .A2(_07924_),
    .B1(net1758),
    .X(_04815_));
 and2_1 _19828_ (.A(_07854_),
    .B(_07921_),
    .X(_04816_));
 or4b_1 _19829_ (.A(_07924_),
    .B(_07925_),
    .C(_04816_),
    .D_N(_07927_),
    .X(_04817_));
 mux2_1 _19830_ (.A0(\digitop_pav2.memctrl_inst.addr_to_reram[2] ),
    .A1(net1759),
    .S(_07931_),
    .X(_01042_));
 mux2_1 _19831_ (.A0(net1140),
    .A1(net1775),
    .S(_07931_),
    .X(_01043_));
 mux2_1 _19832_ (.A0(net1138),
    .A1(_07882_),
    .S(_07931_),
    .X(_01044_));
 and2b_1 _19833_ (.A_N(\digitop_pav2.pie_inst.fsm.past_ctr[7] ),
    .B(\digitop_pav2.pie_inst.fsm.neg_i[7] ),
    .X(_04818_));
 and2b_1 _19834_ (.A_N(\digitop_pav2.pie_inst.fsm.past_ctr[8] ),
    .B(\digitop_pav2.pie_inst.fsm.neg_i[8] ),
    .X(_04819_));
 and2b_1 _19835_ (.A_N(\digitop_pav2.pie_inst.fsm.neg_i[8] ),
    .B(\digitop_pav2.pie_inst.fsm.past_ctr[8] ),
    .X(_04820_));
 nor2_1 _19836_ (.A(_04819_),
    .B(_04820_),
    .Y(_04821_));
 nand2_1 _19837_ (.A(_04818_),
    .B(_04821_),
    .Y(_04822_));
 xnor2_1 _19838_ (.A(_04818_),
    .B(_04821_),
    .Y(_04823_));
 and2b_1 _19839_ (.A_N(\digitop_pav2.pie_inst.fsm.past_ctr[6] ),
    .B(\digitop_pav2.pie_inst.fsm.neg_i[6] ),
    .X(_04824_));
 nand2b_1 _19840_ (.A_N(\digitop_pav2.pie_inst.fsm.past_ctr[6] ),
    .B(\digitop_pav2.pie_inst.fsm.neg_i[6] ),
    .Y(_04825_));
 and2b_1 _19841_ (.A_N(\digitop_pav2.pie_inst.fsm.neg_i[7] ),
    .B(\digitop_pav2.pie_inst.fsm.past_ctr[7] ),
    .X(_04826_));
 or2_1 _19842_ (.A(_04818_),
    .B(_04826_),
    .X(_04827_));
 and2_1 _19843_ (.A(_04825_),
    .B(_04827_),
    .X(_04828_));
 and2b_1 _19844_ (.A_N(\digitop_pav2.pie_inst.fsm.neg_i[6] ),
    .B(\digitop_pav2.pie_inst.fsm.past_ctr[6] ),
    .X(_04829_));
 nor2_1 _19845_ (.A(_04824_),
    .B(_04829_),
    .Y(_04830_));
 and2b_1 _19846_ (.A_N(\digitop_pav2.pie_inst.fsm.past_ctr[5] ),
    .B(\digitop_pav2.pie_inst.fsm.neg_i[5] ),
    .X(_04831_));
 xnor2_1 _19847_ (.A(_04830_),
    .B(_04831_),
    .Y(_04832_));
 and2b_1 _19848_ (.A_N(\digitop_pav2.pie_inst.fsm.past_ctr[4] ),
    .B(\digitop_pav2.pie_inst.fsm.neg_i[4] ),
    .X(_04833_));
 and2b_1 _19849_ (.A_N(\digitop_pav2.pie_inst.fsm.neg_i[5] ),
    .B(\digitop_pav2.pie_inst.fsm.past_ctr[5] ),
    .X(_04834_));
 nor2_1 _19850_ (.A(_04831_),
    .B(_04834_),
    .Y(_04835_));
 nand2_1 _19851_ (.A(_04833_),
    .B(_04835_),
    .Y(_04836_));
 or2_1 _19852_ (.A(_04833_),
    .B(_04835_),
    .X(_04837_));
 nand2_1 _19853_ (.A(_04836_),
    .B(_04837_),
    .Y(_04838_));
 and2b_1 _19854_ (.A_N(\digitop_pav2.pie_inst.fsm.neg_i[4] ),
    .B(\digitop_pav2.pie_inst.fsm.past_ctr[4] ),
    .X(_04839_));
 or4b_1 _19855_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[3] ),
    .B(_04833_),
    .C(_04839_),
    .D_N(\digitop_pav2.pie_inst.fsm.neg_i[3] ),
    .X(_04840_));
 a2bb2o_1 _19856_ (.A1_N(_04833_),
    .A2_N(_04839_),
    .B1(_07148_),
    .B2(\digitop_pav2.pie_inst.fsm.neg_i[3] ),
    .X(_04841_));
 and2_1 _19857_ (.A(_04840_),
    .B(_04841_),
    .X(_04842_));
 xnor2_1 _19858_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[3] ),
    .B(\digitop_pav2.pie_inst.fsm.neg_i[3] ),
    .Y(_04843_));
 and2b_1 _19859_ (.A_N(\digitop_pav2.pie_inst.fsm.past_ctr[2] ),
    .B(\digitop_pav2.pie_inst.fsm.neg_i[2] ),
    .X(_04844_));
 and2b_1 _19860_ (.A_N(\digitop_pav2.pie_inst.fsm.neg_i[2] ),
    .B(\digitop_pav2.pie_inst.fsm.past_ctr[2] ),
    .X(_04845_));
 a211oi_1 _19861_ (.A1(\digitop_pav2.pie_inst.fsm.past_ctr[1] ),
    .A2(_07165_),
    .B1(_04844_),
    .C1(_04845_),
    .Y(_04846_));
 o21a_1 _19862_ (.A1(_04844_),
    .A2(_04846_),
    .B1(_04843_),
    .X(_04847_));
 nand2_1 _19863_ (.A(_04842_),
    .B(_04847_),
    .Y(_04848_));
 a21o_1 _19864_ (.A1(_04840_),
    .A2(_04848_),
    .B1(_04838_),
    .X(_04849_));
 a21oi_1 _19865_ (.A1(_04836_),
    .A2(_04849_),
    .B1(_04832_),
    .Y(_04850_));
 nor2_1 _19866_ (.A(_04825_),
    .B(_04827_),
    .Y(_04851_));
 a211oi_1 _19867_ (.A1(_04830_),
    .A2(_04831_),
    .B1(_04850_),
    .C1(_04851_),
    .Y(_04852_));
 or3_1 _19868_ (.A(_04823_),
    .B(_04828_),
    .C(_04852_),
    .X(_04853_));
 xor2_1 _19869_ (.A(\digitop_pav2.pie_inst.fsm.past_ctr[9] ),
    .B(\digitop_pav2.pie_inst.fsm.neg_i[9] ),
    .X(_04854_));
 xnor2_1 _19870_ (.A(_04819_),
    .B(_04854_),
    .Y(_04855_));
 o21ai_1 _19871_ (.A1(_04828_),
    .A2(_04852_),
    .B1(_04823_),
    .Y(_04856_));
 and3_1 _19872_ (.A(_04832_),
    .B(_04836_),
    .C(_04849_),
    .X(_04857_));
 nor2_1 _19873_ (.A(_04850_),
    .B(_04857_),
    .Y(_04858_));
 xnor2_1 _19874_ (.A(_04842_),
    .B(_04847_),
    .Y(_04859_));
 xnor2_1 _19875_ (.A(_04843_),
    .B(_04844_),
    .Y(_04860_));
 o22a_1 _19876_ (.A1(\digitop_pav2.pie_inst.fsm.past_ctr[1] ),
    .A2(_07165_),
    .B1(_04844_),
    .B2(_04845_),
    .X(_04861_));
 o31a_1 _19877_ (.A1(_04846_),
    .A2(_04860_),
    .A3(_04861_),
    .B1(_04859_),
    .X(_04862_));
 nand3_1 _19878_ (.A(_04838_),
    .B(_04840_),
    .C(_04848_),
    .Y(_04863_));
 nand2_1 _19879_ (.A(_04849_),
    .B(_04863_),
    .Y(_04864_));
 nor2_1 _19880_ (.A(_04862_),
    .B(_04864_),
    .Y(_04865_));
 xor2_1 _19881_ (.A(_04827_),
    .B(_04829_),
    .X(_04866_));
 a21o_1 _19882_ (.A1(_04862_),
    .A2(_04864_),
    .B1(_04866_),
    .X(_04867_));
 a2111o_1 _19883_ (.A1(_04853_),
    .A2(_04856_),
    .B1(_04858_),
    .C1(_04865_),
    .D1(_04867_),
    .X(_04868_));
 a21oi_1 _19884_ (.A1(_04822_),
    .A2(_04853_),
    .B1(_04855_),
    .Y(_04869_));
 a311oi_1 _19885_ (.A1(_04822_),
    .A2(_04853_),
    .A3(_04855_),
    .B1(_04868_),
    .C1(_04869_),
    .Y(_01045_));
 xor2_1 _19886_ (.A(net1103),
    .B(\digitop_pav2.stadly_memctrl_wr_dt9_1.Y ),
    .X(_04870_));
 or2_1 _19887_ (.A(net1099),
    .B(\digitop_pav2.stadly_memctrl_wr_dt10_1.Y ),
    .X(_04871_));
 nand2_1 _19888_ (.A(net1099),
    .B(\digitop_pav2.stadly_memctrl_wr_dt10_1.Y ),
    .Y(_04872_));
 nand2_1 _19889_ (.A(net1087),
    .B(\digitop_pav2.stadly_memctrl_wr_dt14_1.Y ),
    .Y(_04873_));
 or2_1 _19890_ (.A(net1087),
    .B(\digitop_pav2.stadly_memctrl_wr_dt14_1.Y ),
    .X(_04874_));
 nand2_1 _19891_ (.A(net1090),
    .B(\digitop_pav2.stadly_memctrl_wr_dt13_1.Y ),
    .Y(_04875_));
 or2_1 _19892_ (.A(net1090),
    .B(\digitop_pav2.stadly_memctrl_wr_dt13_1.Y ),
    .X(_04876_));
 xor2_1 _19893_ (.A(net1134),
    .B(\digitop_pav2.stadly_memctrl_wr_dt0_1.Y ),
    .X(_04877_));
 nand2_1 _19894_ (.A(net1083),
    .B(\digitop_pav2.stadly_memctrl_wr_dt15_1.Y ),
    .Y(_04878_));
 or2_1 _19895_ (.A(net1083),
    .B(\digitop_pav2.stadly_memctrl_wr_dt15_1.Y ),
    .X(_04879_));
 xor2_1 _19896_ (.A(net1094),
    .B(\digitop_pav2.stadly_memctrl_wr_dt12_1.Y ),
    .X(_04880_));
 a221o_1 _19897_ (.A1(net1131),
    .A2(_07142_),
    .B1(\digitop_pav2.stadly_memctrl_wr_dt2_1.Y ),
    .B2(_07075_),
    .C1(_04880_),
    .X(_04881_));
 xor2_1 _19898_ (.A(net1124),
    .B(\digitop_pav2.stadly_memctrl_wr_dt3_1.Y ),
    .X(_04882_));
 or2_1 _19899_ (.A(net1107),
    .B(\digitop_pav2.stadly_memctrl_wr_dt8_1.Y ),
    .X(_04883_));
 nand2_1 _19900_ (.A(net1107),
    .B(\digitop_pav2.stadly_memctrl_wr_dt8_1.Y ),
    .Y(_04884_));
 o2bb2a_1 _19901_ (.A1_N(_07077_),
    .A2_N(\digitop_pav2.stadly_memctrl_wr_dt5_1.Y ),
    .B1(\digitop_pav2.stadly_memctrl_wr_dt4_1.Y ),
    .B2(_07076_),
    .X(_04885_));
 xor2_1 _19902_ (.A(net1112),
    .B(\digitop_pav2.stadly_memctrl_wr_dt7_1.Y ),
    .X(_04886_));
 a221o_1 _19903_ (.A1(_07076_),
    .A2(\digitop_pav2.stadly_memctrl_wr_dt4_1.Y ),
    .B1(\digitop_pav2.stadly_memctrl_wr_dt6_1.Y ),
    .B2(_07078_),
    .C1(_04870_),
    .X(_04887_));
 or2_1 _19904_ (.A(net1096),
    .B(\digitop_pav2.stadly_memctrl_wr_dt11_1.Y ),
    .X(_04888_));
 nand2_1 _19905_ (.A(net1096),
    .B(\digitop_pav2.stadly_memctrl_wr_dt11_1.Y ),
    .Y(_04889_));
 a221o_1 _19906_ (.A1(net1127),
    .A2(_07143_),
    .B1(_07144_),
    .B2(net1115),
    .C1(_04887_),
    .X(_04890_));
 o221ai_1 _19907_ (.A1(net1131),
    .A2(_07142_),
    .B1(\digitop_pav2.stadly_memctrl_wr_dt5_1.Y ),
    .B2(_07077_),
    .C1(_04885_),
    .Y(_04891_));
 a221o_1 _19908_ (.A1(_04871_),
    .A2(_04872_),
    .B1(_04878_),
    .B2(_04879_),
    .C1(_04886_),
    .X(_04892_));
 a221o_1 _19909_ (.A1(_04883_),
    .A2(_04884_),
    .B1(_04888_),
    .B2(_04889_),
    .C1(_04892_),
    .X(_04893_));
 a211o_1 _19910_ (.A1(_04873_),
    .A2(_04874_),
    .B1(_04891_),
    .C1(_04893_),
    .X(_04894_));
 a211o_1 _19911_ (.A1(_04875_),
    .A2(_04876_),
    .B1(_04890_),
    .C1(_04894_),
    .X(_04895_));
 o41a_2 _19912_ (.A1(_04877_),
    .A2(_04881_),
    .A3(_04882_),
    .A4(_04895_),
    .B1(_07930_),
    .X(_04896_));
 inv_2 _19913_ (.A(_04896_),
    .Y(_04897_));
 nor2_1 _19914_ (.A(_00081_),
    .B(_00079_),
    .Y(_04898_));
 nor2_1 _19915_ (.A(_00081_),
    .B(_00080_),
    .Y(_04899_));
 nor2_1 _19916_ (.A(\digitop_pav2.memctrl_inst.n_state[2] ),
    .B(_04899_),
    .Y(_04900_));
 o21a_1 _19917_ (.A1(_00081_),
    .A2(_00079_),
    .B1(_04900_),
    .X(_04901_));
 and2_1 _19918_ (.A(\digitop_pav2.memctrl_inst.state[1] ),
    .B(_04901_),
    .X(_04902_));
 nand2_1 _19919_ (.A(\digitop_pav2.memctrl_inst.state[1] ),
    .B(_04901_),
    .Y(_04903_));
 nand2_1 _19920_ (.A(net147),
    .B(net145),
    .Y(_04904_));
 or4b_1 _19921_ (.A(\digitop_pav2.memctrl_inst.ctr[7] ),
    .B(\digitop_pav2.memctrl_inst.ctr[6] ),
    .C(_07139_),
    .D_N(\digitop_pav2.memctrl_inst.state[3] ),
    .X(_04905_));
 or4b_4 _19922_ (.A(\digitop_pav2.memctrl_inst.ctr[1] ),
    .B(_09568_),
    .C(_04905_),
    .D_N(\digitop_pav2.memctrl_inst.ctr[0] ),
    .X(_04906_));
 inv_2 _19923_ (.A(_04906_),
    .Y(_04907_));
 or3_1 _19924_ (.A(_07957_),
    .B(_04904_),
    .C(net915),
    .X(_04908_));
 inv_2 _19925_ (.A(net143),
    .Y(_04909_));
 o21a_1 _19926_ (.A1(net1140),
    .A2(_03773_),
    .B1(net1138),
    .X(_04910_));
 nor2_1 _19927_ (.A(net1141),
    .B(net1136),
    .Y(_04911_));
 a22o_1 _19928_ (.A1(net1140),
    .A2(_03790_),
    .B1(net1021),
    .B2(_03781_),
    .X(_04912_));
 o221a_1 _19929_ (.A1(net1026),
    .A2(_03800_),
    .B1(_04910_),
    .B2(_04912_),
    .C1(net914),
    .X(_04913_));
 a31oi_1 _19930_ (.A1(\digitop_pav2.memctrl_inst.flops_0x081[0] ),
    .A2(net149),
    .A3(_04906_),
    .B1(_04913_),
    .Y(_04914_));
 o2bb2a_1 _19931_ (.A1_N(\digitop_pav2.stadly_memctrl_wr_dt0_1.Y ),
    .A2_N(_04896_),
    .B1(net143),
    .B2(_07073_),
    .X(_04915_));
 o21ai_1 _19932_ (.A1(_04904_),
    .A2(_04914_),
    .B1(_04915_),
    .Y(_01047_));
 a22o_1 _19933_ (.A1(net1137),
    .A2(_03825_),
    .B1(net1020),
    .B2(_03809_),
    .X(_04916_));
 a211o_1 _19934_ (.A1(net1140),
    .A2(_03817_),
    .B1(_04916_),
    .C1(_09384_),
    .X(_04917_));
 o211a_1 _19935_ (.A1(net1026),
    .A2(_03837_),
    .B1(net914),
    .C1(_04917_),
    .X(_04918_));
 a31o_1 _19936_ (.A1(\digitop_pav2.memctrl_inst.flops_0x081[1] ),
    .A2(net149),
    .A3(_04906_),
    .B1(_04918_),
    .X(_04919_));
 mux2_1 _19937_ (.A0(net1134),
    .A1(_04919_),
    .S(net145),
    .X(_04920_));
 mux2_1 _19938_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt1_1.Y ),
    .A1(_04920_),
    .S(net147),
    .X(_04921_));
 a21o_1 _19939_ (.A1(net1131),
    .A2(_04909_),
    .B1(_04921_),
    .X(_01048_));
 and3b_1 _19940_ (.A_N(net1141),
    .B(net1138),
    .C(_03856_),
    .X(_04922_));
 a221o_1 _19941_ (.A1(net1141),
    .A2(_03864_),
    .B1(net1020),
    .B2(_03848_),
    .C1(_04922_),
    .X(_04923_));
 nand2_1 _19942_ (.A(_07074_),
    .B(net149),
    .Y(_04924_));
 mux2_1 _19943_ (.A0(_03874_),
    .A1(_04923_),
    .S(net1026),
    .X(_04925_));
 mux2_1 _19944_ (.A0(_04924_),
    .A1(_04925_),
    .S(net914),
    .X(_04926_));
 mux2_1 _19945_ (.A0(net1131),
    .A1(_04926_),
    .S(net146),
    .X(_04927_));
 or2_1 _19946_ (.A(_04896_),
    .B(_04927_),
    .X(_04928_));
 o221a_1 _19947_ (.A1(\digitop_pav2.stadly_memctrl_wr_dt2_1.Y ),
    .A2(net147),
    .B1(net143),
    .B2(net1127),
    .C1(_04928_),
    .X(_01049_));
 a22o_1 _19948_ (.A1(net1139),
    .A2(_03892_),
    .B1(net1021),
    .B2(_03884_),
    .X(_04929_));
 a211o_1 _19949_ (.A1(net1138),
    .A2(_03900_),
    .B1(_04929_),
    .C1(_09384_),
    .X(_04930_));
 and3b_1 _19950_ (.A_N(net149),
    .B(_04906_),
    .C(net67),
    .X(_04931_));
 o211a_1 _19951_ (.A1(net1026),
    .A2(_03910_),
    .B1(net914),
    .C1(_04930_),
    .X(_04932_));
 a31o_1 _19952_ (.A1(\digitop_pav2.memctrl_inst.flops_0x081[3] ),
    .A2(net149),
    .A3(_04906_),
    .B1(_04932_),
    .X(_04933_));
 or3_1 _19953_ (.A(_04902_),
    .B(_04931_),
    .C(_04933_),
    .X(_04934_));
 o211a_1 _19954_ (.A1(net1127),
    .A2(net145),
    .B1(_04934_),
    .C1(net147),
    .X(_04935_));
 a21o_1 _19955_ (.A1(\digitop_pav2.stadly_memctrl_wr_dt3_1.Y ),
    .A2(_04896_),
    .B1(_04909_),
    .X(_04936_));
 o22a_1 _19956_ (.A1(net1124),
    .A2(net143),
    .B1(_04935_),
    .B2(_04936_),
    .X(_01050_));
 a22o_1 _19957_ (.A1(net1137),
    .A2(_03936_),
    .B1(net1020),
    .B2(_03920_),
    .X(_04937_));
 mux2_1 _19958_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.sl_i ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[4] ),
    .S(net150),
    .X(_04938_));
 o21a_1 _19959_ (.A1(net1137),
    .A2(_03928_),
    .B1(net1140),
    .X(_04939_));
 o221a_1 _19960_ (.A1(net1026),
    .A2(_03946_),
    .B1(_04937_),
    .B2(_04939_),
    .C1(net914),
    .X(_04940_));
 a21o_1 _19961_ (.A1(_04906_),
    .A2(_04938_),
    .B1(_04940_),
    .X(_04941_));
 or3_1 _19962_ (.A(net1124),
    .B(_04896_),
    .C(net145),
    .X(_04942_));
 o221a_1 _19963_ (.A1(\digitop_pav2.stadly_memctrl_wr_dt4_1.Y ),
    .A2(net147),
    .B1(_04904_),
    .B2(_04941_),
    .C1(_04942_),
    .X(_04943_));
 mux2_1 _19964_ (.A0(net1122),
    .A1(_04943_),
    .S(net144),
    .X(_01051_));
 mux2_1 _19965_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[5] ),
    .S(net149),
    .X(_04944_));
 and3b_1 _19966_ (.A_N(net1139),
    .B(net1138),
    .C(_03956_),
    .X(_04945_));
 a221o_1 _19967_ (.A1(net1139),
    .A2(_03972_),
    .B1(net1021),
    .B2(_03964_),
    .C1(_04945_),
    .X(_04946_));
 and4b_1 _19968_ (.A_N(net1138),
    .B(net1140),
    .C(\digitop_pav2.memctrl_inst.addr_to_reram[2] ),
    .D(\digitop_pav2.memctrl_inst.addr_to_reram[0] ),
    .X(_04947_));
 mux2_1 _19969_ (.A0(_03982_),
    .A1(_04946_),
    .S(net1026),
    .X(_04948_));
 a211o_1 _19970_ (.A1(\digitop_pav2.memctrl_inst.addr_to_reram[1] ),
    .A2(_04947_),
    .B1(_04948_),
    .C1(_04906_),
    .X(_04949_));
 o21a_1 _19971_ (.A1(net915),
    .A2(_04944_),
    .B1(_04949_),
    .X(_04950_));
 mux2_1 _19972_ (.A0(net1121),
    .A1(_04950_),
    .S(net146),
    .X(_04951_));
 mux2_1 _19973_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt5_1.Y ),
    .A1(_04951_),
    .S(net147),
    .X(_04952_));
 mux2_1 _19974_ (.A0(net1118),
    .A1(_04952_),
    .S(net143),
    .X(_01052_));
 mux2_1 _19975_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_i ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[6] ),
    .S(net150),
    .X(_04953_));
 o21a_1 _19976_ (.A1(net1141),
    .A2(_04000_),
    .B1(net1137),
    .X(_04954_));
 a22o_1 _19977_ (.A1(net1140),
    .A2(_04008_),
    .B1(net1021),
    .B2(_03992_),
    .X(_04955_));
 o2bb2a_1 _19978_ (.A1_N(_09384_),
    .A2_N(_04019_),
    .B1(_04954_),
    .B2(_04955_),
    .X(_04956_));
 mux2_1 _19979_ (.A0(_04953_),
    .A1(_04956_),
    .S(net915),
    .X(_04957_));
 mux2_1 _19980_ (.A0(net1119),
    .A1(_04957_),
    .S(net146),
    .X(_04958_));
 mux2_1 _19981_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt6_1.Y ),
    .A1(_04958_),
    .S(net148),
    .X(_04959_));
 mux2_1 _19982_ (.A0(net1115),
    .A1(_04959_),
    .S(net143),
    .X(_01053_));
 a22o_1 _19983_ (.A1(net1139),
    .A2(_04037_),
    .B1(net1020),
    .B2(_04029_),
    .X(_04960_));
 mux2_1 _19984_ (.A0(\digitop_pav2.invent_inst.s1_i ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[7] ),
    .S(net150),
    .X(_04961_));
 o21a_1 _19985_ (.A1(net1139),
    .A2(_04045_),
    .B1(net1136),
    .X(_04962_));
 o22a_1 _19986_ (.A1(net1026),
    .A2(_04055_),
    .B1(_04960_),
    .B2(_04962_),
    .X(_04963_));
 mux2_1 _19987_ (.A0(_04961_),
    .A1(_04963_),
    .S(net915),
    .X(_04964_));
 mux2_1 _19988_ (.A0(net1115),
    .A1(_04964_),
    .S(net146),
    .X(_04965_));
 mux2_1 _19989_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt7_1.Y ),
    .A1(_04965_),
    .S(net148),
    .X(_04966_));
 mux2_1 _19990_ (.A0(net1111),
    .A1(_04966_),
    .S(net144),
    .X(_01054_));
 a22o_1 _19991_ (.A1(net1139),
    .A2(_04081_),
    .B1(net1021),
    .B2(_04065_),
    .X(_04967_));
 mux2_1 _19992_ (.A0(tclk_i),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[8] ),
    .S(net149),
    .X(_04968_));
 o21a_1 _19993_ (.A1(net1139),
    .A2(_04073_),
    .B1(net1136),
    .X(_04969_));
 o22a_1 _19994_ (.A1(net1026),
    .A2(_04091_),
    .B1(_04967_),
    .B2(_04969_),
    .X(_04970_));
 mux2_1 _19995_ (.A0(_04968_),
    .A1(_04970_),
    .S(net914),
    .X(_04971_));
 mux2_1 _19996_ (.A0(net1111),
    .A1(_04971_),
    .S(net146),
    .X(_04972_));
 mux2_1 _19997_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt8_1.Y ),
    .A1(_04972_),
    .S(net148),
    .X(_04973_));
 mux2_1 _19998_ (.A0(net1107),
    .A1(_04973_),
    .S(net143),
    .X(_01055_));
 a22o_1 _19999_ (.A1(net1137),
    .A2(_04109_),
    .B1(_04117_),
    .B2(net1141),
    .X(_04974_));
 a211o_1 _20000_ (.A1(_04101_),
    .A2(net1020),
    .B1(_04974_),
    .C1(_09384_),
    .X(_04975_));
 and3_1 _20001_ (.A(\digitop_pav2.memctrl_inst.flops_0x081[9] ),
    .B(net149),
    .C(_04906_),
    .X(_04976_));
 o211a_1 _20002_ (.A1(net1026),
    .A2(_04127_),
    .B1(net914),
    .C1(_04975_),
    .X(_04977_));
 o31a_1 _20003_ (.A1(_04931_),
    .A2(_04976_),
    .A3(_04977_),
    .B1(net145),
    .X(_04978_));
 a211o_1 _20004_ (.A1(net1107),
    .A2(_04902_),
    .B1(_04978_),
    .C1(_04896_),
    .X(_04979_));
 o211a_1 _20005_ (.A1(\digitop_pav2.stadly_memctrl_wr_dt9_1.Y ),
    .A2(net147),
    .B1(net143),
    .C1(_04979_),
    .X(_04980_));
 a21o_1 _20006_ (.A1(net1103),
    .A2(_04909_),
    .B1(_04980_),
    .X(_01056_));
 mux2_1 _20007_ (.A0(net1503),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[10] ),
    .S(net150),
    .X(_04981_));
 a22o_1 _20008_ (.A1(net1136),
    .A2(_04145_),
    .B1(_04153_),
    .B2(net1139),
    .X(_04982_));
 a21o_1 _20009_ (.A1(_04137_),
    .A2(net1020),
    .B1(_09384_),
    .X(_04983_));
 o22a_1 _20010_ (.A1(net1027),
    .A2(_04163_),
    .B1(_04982_),
    .B2(_04983_),
    .X(_04984_));
 mux2_1 _20011_ (.A0(_04981_),
    .A1(_04984_),
    .S(net914),
    .X(_04985_));
 mux2_1 _20012_ (.A0(net1104),
    .A1(_04985_),
    .S(net146),
    .X(_04986_));
 mux2_1 _20013_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt10_1.Y ),
    .A1(_04986_),
    .S(net147),
    .X(_04987_));
 mux2_1 _20014_ (.A0(net1099),
    .A1(_04987_),
    .S(net144),
    .X(_01057_));
 a22o_1 _20015_ (.A1(net1139),
    .A2(_04181_),
    .B1(net1020),
    .B2(_04173_),
    .X(_04988_));
 nand2b_1 _20016_ (.A_N(\digitop_pav2.memctrl_inst.flops_0x081[11] ),
    .B(net149),
    .Y(_04989_));
 a211o_1 _20017_ (.A1(net1136),
    .A2(_04189_),
    .B1(_04988_),
    .C1(_09384_),
    .X(_04990_));
 o211a_1 _20018_ (.A1(net1027),
    .A2(_04199_),
    .B1(net914),
    .C1(_04990_),
    .X(_04991_));
 a21oi_1 _20019_ (.A1(_04906_),
    .A2(_04989_),
    .B1(_04991_),
    .Y(_04992_));
 nor2_1 _20020_ (.A(_04902_),
    .B(_04992_),
    .Y(_04993_));
 a211o_1 _20021_ (.A1(net1099),
    .A2(_04902_),
    .B1(_04993_),
    .C1(_04896_),
    .X(_04994_));
 o221a_1 _20022_ (.A1(\digitop_pav2.stadly_memctrl_wr_dt11_1.Y ),
    .A2(net147),
    .B1(net143),
    .B2(net1096),
    .C1(_04994_),
    .X(_01058_));
 mux2_1 _20023_ (.A0(net1746),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[12] ),
    .S(net150),
    .X(_04995_));
 a22o_1 _20024_ (.A1(net1137),
    .A2(_04217_),
    .B1(net1021),
    .B2(_04209_),
    .X(_04996_));
 o21a_1 _20025_ (.A1(net1137),
    .A2(_04225_),
    .B1(net1140),
    .X(_04997_));
 o22a_1 _20026_ (.A1(net1026),
    .A2(_04235_),
    .B1(_04996_),
    .B2(_04997_),
    .X(_04998_));
 mux2_1 _20027_ (.A0(net1747),
    .A1(_04998_),
    .S(net915),
    .X(_04999_));
 mux2_1 _20028_ (.A0(net1096),
    .A1(_04999_),
    .S(net146),
    .X(_05000_));
 mux2_1 _20029_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt12_1.Y ),
    .A1(_05000_),
    .S(net148),
    .X(_05001_));
 mux2_1 _20030_ (.A0(net1094),
    .A1(net1748),
    .S(net144),
    .X(_01059_));
 a22o_1 _20031_ (.A1(net1136),
    .A2(_04253_),
    .B1(net1020),
    .B2(_04245_),
    .X(_05002_));
 mux2_1 _20032_ (.A0(net1738),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[13] ),
    .S(net150),
    .X(_05003_));
 o21a_1 _20033_ (.A1(net1136),
    .A2(_04261_),
    .B1(net1140),
    .X(_05004_));
 o221a_1 _20034_ (.A1(net1027),
    .A2(_04271_),
    .B1(_05002_),
    .B2(_05004_),
    .C1(net914),
    .X(_05005_));
 a21o_1 _20035_ (.A1(_04906_),
    .A2(net1739),
    .B1(_05005_),
    .X(_05006_));
 or3_1 _20036_ (.A(net1094),
    .B(_04896_),
    .C(net145),
    .X(_05007_));
 o221a_1 _20037_ (.A1(\digitop_pav2.stadly_memctrl_wr_dt13_1.Y ),
    .A2(net147),
    .B1(_04904_),
    .B2(_05006_),
    .C1(_05007_),
    .X(_05008_));
 mux2_1 _20038_ (.A0(net1091),
    .A1(net1740),
    .S(net143),
    .X(_01060_));
 mux2_1 _20039_ (.A0(net1743),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[14] ),
    .S(net150),
    .X(_05009_));
 a22o_1 _20040_ (.A1(net1137),
    .A2(_04289_),
    .B1(net1020),
    .B2(_04281_),
    .X(_05010_));
 o21a_1 _20041_ (.A1(net1137),
    .A2(_04297_),
    .B1(net1140),
    .X(_05011_));
 o2bb2a_1 _20042_ (.A1_N(_09384_),
    .A2_N(_04308_),
    .B1(_05010_),
    .B2(_05011_),
    .X(_05012_));
 mux2_1 _20043_ (.A0(net1744),
    .A1(_05012_),
    .S(net915),
    .X(_05013_));
 mux2_1 _20044_ (.A0(net1091),
    .A1(_05013_),
    .S(net146),
    .X(_05014_));
 mux2_1 _20045_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt14_1.Y ),
    .A1(_05014_),
    .S(net148),
    .X(_05015_));
 mux2_1 _20046_ (.A0(net1087),
    .A1(net1745),
    .S(net144),
    .X(_01061_));
 mux2_1 _20047_ (.A0(net1749),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[15] ),
    .S(net150),
    .X(_05016_));
 a22o_1 _20048_ (.A1(net1136),
    .A2(_04326_),
    .B1(net1020),
    .B2(_04318_),
    .X(_05017_));
 o21a_1 _20049_ (.A1(net1136),
    .A2(_04334_),
    .B1(net1141),
    .X(_05018_));
 o2bb2a_1 _20050_ (.A1_N(_09384_),
    .A2_N(_04345_),
    .B1(_05017_),
    .B2(_05018_),
    .X(_05019_));
 mux2_1 _20051_ (.A0(_05016_),
    .A1(_05019_),
    .S(net915),
    .X(_05020_));
 mux2_1 _20052_ (.A0(net1087),
    .A1(_05020_),
    .S(net146),
    .X(_05021_));
 mux2_1 _20053_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt15_1.Y ),
    .A1(_05021_),
    .S(net148),
    .X(_05022_));
 mux2_1 _20054_ (.A0(net1084),
    .A1(net1750),
    .S(net144),
    .X(_01062_));
 a21oi_1 _20055_ (.A1(\digitop_pav2.memctrl_inst.bit_addr[0] ),
    .A2(net145),
    .B1(_10320_),
    .Y(_05023_));
 o21ai_1 _20056_ (.A1(\digitop_pav2.memctrl_inst.bit_addr[0] ),
    .A2(net145),
    .B1(_05023_),
    .Y(_01063_));
 o21a_1 _20057_ (.A1(\digitop_pav2.memctrl_inst.bit_addr[0] ),
    .A2(net145),
    .B1(\digitop_pav2.memctrl_inst.bit_addr[1] ),
    .X(_05024_));
 or3_1 _20058_ (.A(\digitop_pav2.memctrl_inst.bit_addr[0] ),
    .B(\digitop_pav2.memctrl_inst.bit_addr[1] ),
    .C(net145),
    .X(_05025_));
 or3b_1 _20059_ (.A(_10320_),
    .B(_05024_),
    .C_N(_05025_),
    .X(_01064_));
 or2_1 _20060_ (.A(\digitop_pav2.memctrl_inst.bit_addr[2] ),
    .B(_05025_),
    .X(_05026_));
 nand2_1 _20061_ (.A(_10321_),
    .B(_05026_),
    .Y(_05027_));
 a21o_1 _20062_ (.A1(\digitop_pav2.memctrl_inst.bit_addr[2] ),
    .A2(_05025_),
    .B1(_05027_),
    .X(_01065_));
 xor2_1 _20063_ (.A(\digitop_pav2.memctrl_inst.bit_addr[3] ),
    .B(_05026_),
    .X(_05028_));
 nand2_1 _20064_ (.A(_10321_),
    .B(_05028_),
    .Y(_01066_));
 and3b_1 _20065_ (.A_N(\digitop_pav2.memctrl_inst.n_state[2] ),
    .B(_00079_),
    .C(_04899_),
    .X(_05029_));
 nand2_1 _20066_ (.A(\digitop_pav2.memctrl_inst.state[2] ),
    .B(_05029_),
    .Y(_05030_));
 a31o_1 _20067_ (.A1(_07139_),
    .A2(_09572_),
    .A3(_05030_),
    .B1(_09571_),
    .X(_05031_));
 and2_1 _20068_ (.A(\digitop_pav2.memctrl_inst.state[0] ),
    .B(_05029_),
    .X(_05032_));
 a31o_1 _20069_ (.A1(\digitop_pav2.memctrl_inst.state[0] ),
    .A2(_04898_),
    .A3(_04900_),
    .B1(_05032_),
    .X(_05033_));
 o21a_1 _20070_ (.A1(\digitop_pav2.memctrl_inst.state[1] ),
    .A2(\digitop_pav2.memctrl_inst.state[2] ),
    .B1(_04901_),
    .X(_05034_));
 inv_2 _20071_ (.A(_05034_),
    .Y(_05035_));
 nor2_1 _20072_ (.A(_05033_),
    .B(_05034_),
    .Y(_05036_));
 and2_1 _20073_ (.A(_05031_),
    .B(_05036_),
    .X(_05037_));
 nand2_1 _20074_ (.A(_05031_),
    .B(_05036_),
    .Y(_05038_));
 a21oi_1 _20075_ (.A1(\digitop_pav2.memctrl_inst.ctr[0] ),
    .A2(_05035_),
    .B1(_05033_),
    .Y(_05039_));
 mux2_1 _20076_ (.A0(\digitop_pav2.memctrl_inst.ctr[0] ),
    .A1(_05039_),
    .S(_05038_),
    .X(_01067_));
 nor2_1 _20077_ (.A(_05032_),
    .B(_05037_),
    .Y(_05040_));
 nand2_1 _20078_ (.A(\digitop_pav2.memctrl_inst.ctr[0] ),
    .B(\digitop_pav2.memctrl_inst.ctr[1] ),
    .Y(_05041_));
 nand3_1 _20079_ (.A(_09566_),
    .B(_05036_),
    .C(_05041_),
    .Y(_05042_));
 a22o_1 _20080_ (.A1(\digitop_pav2.memctrl_inst.ctr[1] ),
    .A2(_05037_),
    .B1(_05040_),
    .B2(_05042_),
    .X(_01068_));
 or2_1 _20081_ (.A(\digitop_pav2.memctrl_inst.ctr[2] ),
    .B(_09566_),
    .X(_05043_));
 nand2_1 _20082_ (.A(\digitop_pav2.memctrl_inst.ctr[2] ),
    .B(_09566_),
    .Y(_05044_));
 a311o_1 _20083_ (.A1(_05035_),
    .A2(_05043_),
    .A3(_05044_),
    .B1(_05037_),
    .C1(_05033_),
    .X(_05045_));
 a21bo_1 _20084_ (.A1(\digitop_pav2.memctrl_inst.ctr[2] ),
    .A2(_05037_),
    .B1_N(_05045_),
    .X(_01069_));
 nor4_1 _20085_ (.A(\digitop_pav2.memctrl_inst.ctr[2] ),
    .B(\digitop_pav2.memctrl_inst.ctr[3] ),
    .C(_09566_),
    .D(_05031_),
    .Y(_05046_));
 o31a_1 _20086_ (.A1(\digitop_pav2.memctrl_inst.ctr[2] ),
    .A2(_09566_),
    .A3(_05031_),
    .B1(\digitop_pav2.memctrl_inst.ctr[3] ),
    .X(_05047_));
 o21a_1 _20087_ (.A1(_05046_),
    .A2(_05047_),
    .B1(_05036_),
    .X(_01070_));
 nand2_1 _20088_ (.A(\digitop_pav2.memctrl_inst.ctr[4] ),
    .B(net142),
    .Y(_05048_));
 o211a_1 _20089_ (.A1(\digitop_pav2.memctrl_inst.ctr[4] ),
    .A2(net142),
    .B1(_05048_),
    .C1(_05036_),
    .X(_01071_));
 o21ai_1 _20090_ (.A1(_09566_),
    .A2(_09567_),
    .B1(\digitop_pav2.memctrl_inst.ctr[5] ),
    .Y(_05049_));
 a211o_1 _20091_ (.A1(_09569_),
    .A2(_05049_),
    .B1(_05034_),
    .C1(_05033_),
    .X(_05050_));
 o2bb2a_1 _20092_ (.A1_N(_05040_),
    .A2_N(_05050_),
    .B1(\digitop_pav2.memctrl_inst.ctr[5] ),
    .B2(_05038_),
    .X(_01072_));
 nand2_1 _20093_ (.A(\digitop_pav2.memctrl_inst.ctr[6] ),
    .B(_09569_),
    .Y(_05051_));
 a211o_1 _20094_ (.A1(_09570_),
    .A2(_05051_),
    .B1(_05034_),
    .C1(_05033_),
    .X(_05052_));
 o2bb2a_1 _20095_ (.A1_N(_05040_),
    .A2_N(_05052_),
    .B1(\digitop_pav2.memctrl_inst.ctr[6] ),
    .B2(_05038_),
    .X(_01073_));
 and2_1 _20096_ (.A(\digitop_pav2.memctrl_inst.ctr[7] ),
    .B(_09570_),
    .X(_05053_));
 o21ai_1 _20097_ (.A1(_09571_),
    .A2(_05053_),
    .B1(_05036_),
    .Y(_05054_));
 o2bb2a_1 _20098_ (.A1_N(_05040_),
    .A2_N(_05054_),
    .B1(\digitop_pav2.memctrl_inst.ctr[7] ),
    .B2(_05038_),
    .X(_01074_));
 o21bai_1 _20099_ (.A1(\digitop_pav2.memctrl_inst.nvm_rd_en_i ),
    .A2(_10321_),
    .B1_N(\digitop_pav2.func_reg_wr_en ),
    .Y(_01075_));
 o21a_1 _20100_ (.A1(\digitop_pav2.memctrl_inst.bit_addr_allow ),
    .A2(_10320_),
    .B1(\digitop_pav2.memctrl_inst.n_bit_addr_allow ),
    .X(_01076_));
 mux2_1 _20101_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[0] ),
    .A1(_08520_),
    .S(net530),
    .X(_01079_));
 mux2_1 _20102_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[0] ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[1] ),
    .S(net531),
    .X(_01080_));
 mux2_1 _20103_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[2] ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[1] ),
    .S(net530),
    .X(_01081_));
 mux2_1 _20104_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[2] ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[3] ),
    .S(net532),
    .X(_01082_));
 mux2_1 _20105_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[3] ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[4] ),
    .S(net532),
    .X(_01083_));
 mux2_1 _20106_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[4] ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[5] ),
    .S(net532),
    .X(_01084_));
 mux2_1 _20107_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[6] ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[5] ),
    .S(_09541_),
    .X(_01085_));
 nor3_1 _20108_ (.A(net1274),
    .B(net1672),
    .C(net1279),
    .Y(_05055_));
 o32a_1 _20109_ (.A1(net1247),
    .A2(net1715),
    .A3(_05055_),
    .B1(_07654_),
    .B2(_07063_),
    .X(_05056_));
 a211o_1 _20110_ (.A1(_00170_),
    .A2(_08982_),
    .B1(_09003_),
    .C1(_08980_),
    .X(_05057_));
 or3b_1 _20111_ (.A(_00170_),
    .B(net974),
    .C_N(_09001_),
    .X(_05058_));
 nand3_1 _20112_ (.A(_08967_),
    .B(_05057_),
    .C(_05058_),
    .Y(_05059_));
 o211a_1 _20113_ (.A1(\digitop_pav2.invent_inst.s1_r_o ),
    .A2(_08967_),
    .B1(_05056_),
    .C1(_05059_),
    .X(_01086_));
 and3b_1 _20114_ (.A_N(net974),
    .B(_09001_),
    .C(_00170_),
    .X(_05060_));
 o221a_1 _20115_ (.A1(\digitop_pav2.invent_inst.s1_s_o ),
    .A2(_08967_),
    .B1(_09006_),
    .B2(_05060_),
    .C1(_05056_),
    .X(_01090_));
 nor2_1 _20116_ (.A(_10339_),
    .B(_03682_),
    .Y(_05061_));
 mux2_1 _20117_ (.A0(net1178),
    .A1(net814),
    .S(_05061_),
    .X(_01093_));
 nor2_1 _20118_ (.A(_10339_),
    .B(_03665_),
    .Y(_05062_));
 mux2_1 _20119_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[7] ),
    .A1(net815),
    .S(_05062_),
    .X(_01094_));
 or2_1 _20120_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[3] ),
    .B(_07135_),
    .X(_05063_));
 nand2_1 _20121_ (.A(net802),
    .B(_05063_),
    .Y(_05064_));
 o22a_1 _20122_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[4] ),
    .A2(_10339_),
    .B1(_03667_),
    .B2(_10333_),
    .X(_05065_));
 nor2_1 _20123_ (.A(_10334_),
    .B(_03666_),
    .Y(_05066_));
 o21ai_1 _20124_ (.A1(_03663_),
    .A2(_05066_),
    .B1(_05065_),
    .Y(_05067_));
 a211o_1 _20125_ (.A1(_07135_),
    .A2(_03674_),
    .B1(_05067_),
    .C1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[3] ),
    .X(_05068_));
 xnor2_1 _20126_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[1] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[2] ),
    .Y(_05069_));
 o22a_1 _20127_ (.A1(_03663_),
    .A2(_03670_),
    .B1(_03674_),
    .B2(_10340_),
    .X(_05070_));
 mux2_1 _20128_ (.A0(_10333_),
    .A1(_05070_),
    .S(_05069_),
    .X(_05071_));
 o211ai_1 _20129_ (.A1(_10340_),
    .A2(_03675_),
    .B1(_05068_),
    .C1(_05071_),
    .Y(_05072_));
 mux2_1 _20130_ (.A0(_05072_),
    .A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[0] ),
    .S(_05064_),
    .X(_01095_));
 a21o_1 _20131_ (.A1(_10333_),
    .A2(_03674_),
    .B1(_10334_),
    .X(_05073_));
 a2bb2o_1 _20132_ (.A1_N(_10333_),
    .A2_N(_03667_),
    .B1(_05063_),
    .B2(_05073_),
    .X(_05074_));
 mux2_1 _20133_ (.A0(_05074_),
    .A1(net1177),
    .S(_05064_),
    .X(_01096_));
 or2_1 _20134_ (.A(net1176),
    .B(_10334_),
    .X(_05075_));
 a31o_1 _20135_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[3] ),
    .A2(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[4] ),
    .A3(_05075_),
    .B1(_05067_),
    .X(_05076_));
 mux2_1 _20136_ (.A0(_05076_),
    .A1(net1176),
    .S(_05064_),
    .X(_01097_));
 o21bai_1 _20137_ (.A1(_05064_),
    .A2(_05065_),
    .B1_N(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[3] ),
    .Y(_01098_));
 a31o_1 _20138_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[3] ),
    .A2(net802),
    .A3(_03672_),
    .B1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[4] ),
    .X(_01099_));
 a31o_1 _20139_ (.A1(net974),
    .A2(_08977_),
    .A3(_09004_),
    .B1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s0_i ),
    .X(_05077_));
 or3_1 _20140_ (.A(_07127_),
    .B(_08968_),
    .C(_08969_),
    .X(_05078_));
 o31a_1 _20141_ (.A1(net1179),
    .A2(net1180),
    .A3(\digitop_pav2.dr ),
    .B1(net1272),
    .X(_05079_));
 a31o_1 _20142_ (.A1(net1272),
    .A2(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[5] ),
    .A3(_10675_),
    .B1(_08978_),
    .X(_05080_));
 o31ai_1 _20143_ (.A1(_07063_),
    .A2(\digitop_pav2.invent_inst.invent_sel_pav2.mask_mismatch_ff ),
    .A3(_08975_),
    .B1(_05080_),
    .Y(_05081_));
 mux2_1 _20144_ (.A0(_05078_),
    .A1(_05079_),
    .S(net974),
    .X(_05082_));
 a21bo_1 _20145_ (.A1(net974),
    .A2(_05081_),
    .B1_N(_05077_),
    .X(_05083_));
 mux2_1 _20146_ (.A0(_05083_),
    .A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.s0_i ),
    .S(_05082_),
    .X(_01100_));
 a21o_1 _20147_ (.A1(_10341_),
    .A2(_10397_),
    .B1(_03684_),
    .X(_05084_));
 and2_1 _20148_ (.A(_04470_),
    .B(_05084_),
    .X(_05085_));
 mux2_1 _20149_ (.A0(_07137_),
    .A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[6] ),
    .S(net1013),
    .X(_05086_));
 mux2_1 _20150_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[0] ),
    .A1(_05086_),
    .S(net526),
    .X(_01101_));
 a21oi_1 _20151_ (.A1(_10408_),
    .A2(_10578_),
    .B1(net1013),
    .Y(_05087_));
 a21o_1 _20152_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[5] ),
    .A2(net1013),
    .B1(_05087_),
    .X(_05088_));
 mux2_1 _20153_ (.A0(net1175),
    .A1(_05088_),
    .S(net526),
    .X(_01102_));
 xor2_1 _20154_ (.A(net1174),
    .B(_10570_),
    .X(_05089_));
 nor2_1 _20155_ (.A(net1012),
    .B(_05089_),
    .Y(_05090_));
 a31o_1 _20156_ (.A1(net1270),
    .A2(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[4] ),
    .A3(net1013),
    .B1(_05090_),
    .X(_05091_));
 mux2_1 _20157_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[2] ),
    .A1(_05091_),
    .S(net526),
    .X(_01103_));
 a31o_1 _20158_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[0] ),
    .A2(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[1] ),
    .A3(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[2] ),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[3] ),
    .X(_05092_));
 nor3b_1 _20159_ (.A(_10571_),
    .B(net1012),
    .C_N(_05092_),
    .Y(_05093_));
 a31o_1 _20160_ (.A1(net1270),
    .A2(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[3] ),
    .A3(net1012),
    .B1(_05093_),
    .X(_05094_));
 mux2_1 _20161_ (.A0(net1173),
    .A1(_05094_),
    .S(_05085_),
    .X(_01104_));
 o21bai_1 _20162_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[4] ),
    .A2(_10571_),
    .B1_N(net1012),
    .Y(_05095_));
 a2bb2o_1 _20163_ (.A1_N(_10634_),
    .A2_N(_05095_),
    .B1(net1012),
    .B2(_07857_),
    .X(_05096_));
 mux2_1 _20164_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[4] ),
    .A1(_05096_),
    .S(net526),
    .X(_01105_));
 or2_1 _20165_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[5] ),
    .B(_10634_),
    .X(_05097_));
 a21oi_1 _20166_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[5] ),
    .A2(_10634_),
    .B1(net1012),
    .Y(_05098_));
 a22o_1 _20167_ (.A1(_07858_),
    .A2(net1012),
    .B1(_05097_),
    .B2(_05098_),
    .X(_05099_));
 mux2_1 _20168_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[5] ),
    .A1(_05099_),
    .S(net526),
    .X(_01106_));
 a31o_1 _20169_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[4] ),
    .A2(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[5] ),
    .A3(_10571_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[6] ),
    .X(_05100_));
 and3_1 _20170_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[5] ),
    .B(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[6] ),
    .C(_10634_),
    .X(_05101_));
 nor2_1 _20171_ (.A(net1012),
    .B(_05101_),
    .Y(_05102_));
 a22o_1 _20172_ (.A1(_07860_),
    .A2(net1012),
    .B1(_05100_),
    .B2(_05102_),
    .X(_05103_));
 mux2_1 _20173_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[6] ),
    .A1(_05103_),
    .S(net526),
    .X(_01107_));
 a21o_1 _20174_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[7] ),
    .A2(_05101_),
    .B1(net1012),
    .X(_05104_));
 a21oi_1 _20175_ (.A1(net526),
    .A2(_05101_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[7] ),
    .Y(_05105_));
 a21oi_1 _20176_ (.A1(net526),
    .A2(_05104_),
    .B1(_05105_),
    .Y(_01108_));
 a21boi_1 _20177_ (.A1(net526),
    .A2(_05104_),
    .B1_N(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[8] ),
    .Y(_05106_));
 nor2_1 _20178_ (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[8] ),
    .B(net1013),
    .Y(_05107_));
 a41o_1 _20179_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[7] ),
    .A2(net526),
    .A3(_05101_),
    .A4(_05107_),
    .B1(_05106_),
    .X(_01109_));
 nand2_1 _20180_ (.A(net159),
    .B(_04472_),
    .Y(_05108_));
 a221oi_1 _20181_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[7] ),
    .A2(_07901_),
    .B1(_07902_),
    .B2(\digitop_pav2.invent_inst.invent_sel_pav2.state[11] ),
    .C1(_05108_),
    .Y(_05109_));
 o211a_1 _20182_ (.A1(_07909_),
    .A2(_04471_),
    .B1(_05109_),
    .C1(_04470_),
    .X(_05110_));
 mux2_1 _20183_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[0] ),
    .A1(net1135),
    .S(net153),
    .X(_01110_));
 mux2_1 _20184_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[1] ),
    .A1(net1133),
    .S(net154),
    .X(_01111_));
 mux2_1 _20185_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[2] ),
    .A1(net1129),
    .S(net153),
    .X(_01112_));
 mux2_1 _20186_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[3] ),
    .A1(net1125),
    .S(net153),
    .X(_01113_));
 mux2_1 _20187_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[4] ),
    .A1(net1122),
    .S(net154),
    .X(_01114_));
 mux2_1 _20188_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[5] ),
    .A1(net1119),
    .S(net153),
    .X(_01115_));
 mux2_1 _20189_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[6] ),
    .A1(net1116),
    .S(net153),
    .X(_01116_));
 mux2_1 _20190_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[7] ),
    .A1(net1113),
    .S(net153),
    .X(_01117_));
 mux2_1 _20191_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[8] ),
    .A1(net1109),
    .S(net153),
    .X(_01118_));
 mux2_1 _20192_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[9] ),
    .A1(net1105),
    .S(net154),
    .X(_01119_));
 mux2_1 _20193_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[10] ),
    .A1(net1101),
    .S(net154),
    .X(_01120_));
 mux2_1 _20194_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[11] ),
    .A1(net1097),
    .S(net154),
    .X(_01121_));
 mux2_1 _20195_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[12] ),
    .A1(net1095),
    .S(net154),
    .X(_01122_));
 mux2_1 _20196_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[13] ),
    .A1(net1092),
    .S(net153),
    .X(_01123_));
 mux2_1 _20197_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[14] ),
    .A1(net1088),
    .S(net153),
    .X(_01124_));
 mux2_1 _20198_ (.A0(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[15] ),
    .A1(net1085),
    .S(net153),
    .X(_01125_));
 o21a_1 _20199_ (.A1(\digitop_pav2.invent_inst.invent_sel_pav2.state[9] ),
    .A2(_10565_),
    .B1(_10325_),
    .X(_05111_));
 a31o_1 _20200_ (.A1(_10648_),
    .A2(net802),
    .A3(_05111_),
    .B1(\digitop_pav2.invent_inst.invent_sel_pav2.mask_mismatch_ff ),
    .X(_01126_));
 or2_1 _20201_ (.A(net1169),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[3] ),
    .X(_05112_));
 or2_1 _20202_ (.A(net1168),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[3] ),
    .X(_05113_));
 or2_1 _20203_ (.A(net1169),
    .B(_05113_),
    .X(_05114_));
 or2_2 _20204_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[0] ),
    .B(_05114_),
    .X(_05115_));
 nor2_1 _20205_ (.A(net1170),
    .B(net1164),
    .Y(_05116_));
 or2_1 _20206_ (.A(net1170),
    .B(net1164),
    .X(_05117_));
 mux2_1 _20207_ (.A0(net1171),
    .A1(net1165),
    .S(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[0] ),
    .X(_05118_));
 a31o_1 _20208_ (.A1(net1737),
    .A2(_05115_),
    .A3(_05116_),
    .B1(_05118_),
    .X(_01127_));
 nand2_1 _20209_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[0] ),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[1] ),
    .Y(_05119_));
 nand2_1 _20210_ (.A(_10682_),
    .B(_05119_),
    .Y(_05120_));
 a22o_1 _20211_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[1] ),
    .A2(net1164),
    .B1(_05120_),
    .B2(net1170),
    .X(_05121_));
 a31o_1 _20212_ (.A1(net1735),
    .A2(_05114_),
    .A3(_05116_),
    .B1(_05121_),
    .X(_01128_));
 and2_2 _20213_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[0] ),
    .B(net1169),
    .X(_05122_));
 o21a_1 _20214_ (.A1(_05113_),
    .A2(_05122_),
    .B1(_08891_),
    .X(_05123_));
 o21ai_1 _20215_ (.A1(net1164),
    .A2(_10682_),
    .B1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[2] ),
    .Y(_05124_));
 o31a_1 _20216_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[2] ),
    .A2(net1164),
    .A3(_10682_),
    .B1(_05117_),
    .X(_05125_));
 o2bb2a_1 _20217_ (.A1_N(_05124_),
    .A2_N(_05125_),
    .B1(_05117_),
    .B2(_05123_),
    .X(_01129_));
 nand2_1 _20218_ (.A(_05113_),
    .B(_05116_),
    .Y(_05126_));
 or4b_1 _20219_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[2] ),
    .B(_10682_),
    .C(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[3] ),
    .D_N(net1170),
    .X(_05127_));
 o21a_1 _20220_ (.A1(net1742),
    .A2(_05126_),
    .B1(_05127_),
    .X(_05128_));
 a21bo_1 _20221_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[3] ),
    .A2(_05125_),
    .B1_N(_05128_),
    .X(_01130_));
 o211a_1 _20222_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[0] ),
    .A2(_05112_),
    .B1(_05113_),
    .C1(_05116_),
    .X(_05129_));
 a2bb2o_1 _20223_ (.A1_N(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[4] ),
    .A2_N(_05127_),
    .B1(_05129_),
    .B2(_08890_),
    .X(_05130_));
 a31o_1 _20224_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[4] ),
    .A2(_05117_),
    .A3(_05127_),
    .B1(_05130_),
    .X(_01131_));
 o21ai_1 _20225_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[5] ),
    .A2(_10683_),
    .B1(net1170),
    .Y(_05131_));
 nand2_1 _20226_ (.A(_07339_),
    .B(_05131_),
    .Y(_05132_));
 a31o_1 _20227_ (.A1(_08895_),
    .A2(_05112_),
    .A3(_05113_),
    .B1(_05117_),
    .X(_05133_));
 a21o_1 _20228_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[5] ),
    .A2(_10683_),
    .B1(_05131_),
    .X(_05134_));
 o211a_1 _20229_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[5] ),
    .A2(_07339_),
    .B1(_05133_),
    .C1(_05134_),
    .X(_01132_));
 o2111a_1 _20230_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[3] ),
    .A2(_05122_),
    .B1(_05116_),
    .C1(_05113_),
    .D1(_08900_),
    .X(_05135_));
 a221o_1 _20231_ (.A1(net1170),
    .A2(_10685_),
    .B1(_05132_),
    .B2(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[6] ),
    .C1(_05135_),
    .X(_01133_));
 xnor2_1 _20232_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[7] ),
    .B(_10684_),
    .Y(_05136_));
 and2b_1 _20233_ (.A_N(net1171),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[3] ),
    .X(_05137_));
 a31o_1 _20234_ (.A1(net1476),
    .A2(net1732),
    .A3(_05137_),
    .B1(net1164),
    .X(_05138_));
 or2_1 _20235_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[7] ),
    .B(_07339_),
    .X(_05139_));
 a22o_1 _20236_ (.A1(net1170),
    .A2(_05136_),
    .B1(net1733),
    .B2(_05139_),
    .X(_01134_));
 o21ai_1 _20237_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[7] ),
    .A2(_10684_),
    .B1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[8] ),
    .Y(_05140_));
 nand2_1 _20238_ (.A(_10686_),
    .B(_05140_),
    .Y(_05141_));
 o31a_1 _20239_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[0] ),
    .A2(net1169),
    .A3(net1168),
    .B1(_05137_),
    .X(_05142_));
 and3_1 _20240_ (.A(_07339_),
    .B(_08903_),
    .C(_05142_),
    .X(_05143_));
 a221o_1 _20241_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[8] ),
    .A2(net1164),
    .B1(_05141_),
    .B2(net1170),
    .C1(_05143_),
    .X(_01135_));
 nand2_1 _20242_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[9] ),
    .B(_10686_),
    .Y(_05144_));
 a21boi_1 _20243_ (.A1(_10687_),
    .A2(_05144_),
    .B1_N(net1170),
    .Y(_05145_));
 o2111a_1 _20244_ (.A1(net1169),
    .A2(net1168),
    .B1(_07339_),
    .C1(_08911_),
    .D1(_05137_),
    .X(_05146_));
 a211o_1 _20245_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[9] ),
    .A2(net1164),
    .B1(_05145_),
    .C1(_05146_),
    .X(_01136_));
 xnor2_1 _20246_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[10] ),
    .B(_10687_),
    .Y(_05147_));
 o2111a_1 _20247_ (.A1(net1168),
    .A2(_05122_),
    .B1(_05137_),
    .C1(_07339_),
    .D1(_08908_),
    .X(_05148_));
 a221o_1 _20248_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[10] ),
    .A2(net1165),
    .B1(_05147_),
    .B2(net1171),
    .C1(_05148_),
    .X(_01137_));
 o21ai_1 _20249_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[10] ),
    .A2(_10687_),
    .B1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[11] ),
    .Y(_05149_));
 nand2_1 _20250_ (.A(_10688_),
    .B(_05149_),
    .Y(_05150_));
 a32o_1 _20251_ (.A1(net1168),
    .A2(_08913_),
    .A3(_05137_),
    .B1(_05150_),
    .B2(net1170),
    .X(_05151_));
 mux2_1 _20252_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[11] ),
    .A1(_05151_),
    .S(_07339_),
    .X(_01138_));
 nand2_1 _20253_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[12] ),
    .B(_10688_),
    .Y(_05152_));
 a21boi_1 _20254_ (.A1(_10689_),
    .A2(_05152_),
    .B1_N(net1171),
    .Y(_05153_));
 and3_1 _20255_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[9] ),
    .B(net1168),
    .C(_05137_),
    .X(_05154_));
 o211a_1 _20256_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[0] ),
    .A2(net1169),
    .B1(_08909_),
    .C1(_05154_),
    .X(_05155_));
 a211o_1 _20257_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[12] ),
    .A2(net1164),
    .B1(_05153_),
    .C1(_05155_),
    .X(_01139_));
 and2_1 _20258_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[13] ),
    .B(_10689_),
    .X(_05156_));
 o21a_1 _20259_ (.A1(_10690_),
    .A2(_05156_),
    .B1(net1171),
    .X(_05157_));
 a41o_1 _20260_ (.A1(net1169),
    .A2(net1168),
    .A3(_08883_),
    .A4(_05137_),
    .B1(net1165),
    .X(_05158_));
 o22a_1 _20261_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[13] ),
    .A2(_07339_),
    .B1(_05157_),
    .B2(_05158_),
    .X(_01140_));
 o21a_1 _20262_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[13] ),
    .A2(_10689_),
    .B1(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[14] ),
    .X(_05159_));
 o21a_1 _20263_ (.A1(_10691_),
    .A2(_05159_),
    .B1(net1171),
    .X(_05160_));
 a32o_1 _20264_ (.A1(_08881_),
    .A2(_05122_),
    .A3(_05154_),
    .B1(net1164),
    .B2(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[14] ),
    .X(_05161_));
 or2_1 _20265_ (.A(_05160_),
    .B(_05161_),
    .X(_01141_));
 nand2_1 _20266_ (.A(_10341_),
    .B(net802),
    .Y(_05162_));
 mux2_1 _20267_ (.A0(net814),
    .A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[7] ),
    .S(_05162_),
    .X(_01142_));
 mux2_1 _20268_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.query_inversion ),
    .A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.flags_en_o ),
    .S(_08999_),
    .X(_01143_));
 a31o_1 _20269_ (.A1(net1168),
    .A2(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[3] ),
    .A3(_05122_),
    .B1(_08975_),
    .X(_05163_));
 nand2_1 _20270_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[4] ),
    .B(_05163_),
    .Y(_05164_));
 a21oi_1 _20271_ (.A1(_08973_),
    .A2(_05115_),
    .B1(_05164_),
    .Y(_05165_));
 o21ba_2 _20272_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[7] ),
    .A2(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[4] ),
    .B1_N(_05165_),
    .X(_05166_));
 inv_2 _20273_ (.A(_05166_),
    .Y(_05167_));
 mux2_1 _20274_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[4] ),
    .A1(_07136_),
    .S(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[4] ),
    .X(_05168_));
 mux2_1 _20275_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[0] ),
    .A1(_05168_),
    .S(_05166_),
    .X(_01144_));
 or2_1 _20276_ (.A(net1169),
    .B(_08973_),
    .X(_05169_));
 nand2_1 _20277_ (.A(net1169),
    .B(_08973_),
    .Y(_05170_));
 a21oi_1 _20278_ (.A1(_05169_),
    .A2(_05170_),
    .B1(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[0] ),
    .Y(_05171_));
 and3_1 _20279_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[0] ),
    .B(_05169_),
    .C(_05170_),
    .X(_05172_));
 nor2_1 _20280_ (.A(_05171_),
    .B(_05172_),
    .Y(_05173_));
 mux2_1 _20281_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[3] ),
    .A1(_05173_),
    .S(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[4] ),
    .X(_05174_));
 mux2_1 _20282_ (.A0(net1169),
    .A1(_05174_),
    .S(_05166_),
    .X(_01145_));
 nor2_1 _20283_ (.A(net1168),
    .B(_08973_),
    .Y(_05175_));
 and3_1 _20284_ (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[3] ),
    .B(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[4] ),
    .C(net1168),
    .X(_05176_));
 nor2_1 _20285_ (.A(_05175_),
    .B(_05176_),
    .Y(_05177_));
 a21o_1 _20286_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[1] ),
    .A2(_08973_),
    .B1(_05172_),
    .X(_05178_));
 xnor2_1 _20287_ (.A(_05177_),
    .B(_05178_),
    .Y(_05179_));
 nand2_1 _20288_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[4] ),
    .B(_05179_),
    .Y(_05180_));
 o21a_1 _20289_ (.A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[2] ),
    .A2(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[4] ),
    .B1(_05166_),
    .X(_05181_));
 a22o_1 _20290_ (.A1(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[2] ),
    .A2(_05167_),
    .B1(_05180_),
    .B2(_05181_),
    .X(_01146_));
 a21oi_1 _20291_ (.A1(_05177_),
    .A2(_05178_),
    .B1(_05176_),
    .Y(_05182_));
 xor2_1 _20292_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[3] ),
    .B(_08973_),
    .X(_05183_));
 xnor2_1 _20293_ (.A(_05182_),
    .B(_05183_),
    .Y(_05184_));
 mux2_1 _20294_ (.A0(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[1] ),
    .A1(_05184_),
    .S(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[4] ),
    .X(_05185_));
 mux2_1 _20295_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[3] ),
    .A1(_05185_),
    .S(_05166_),
    .X(_01147_));
 and2_1 _20296_ (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[7] ),
    .B(_08999_),
    .X(_05186_));
 mux2_1 _20297_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[0] ),
    .A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[7] ),
    .S(_05186_),
    .X(_01148_));
 mux2_1 _20298_ (.A0(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[1] ),
    .A1(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[6] ),
    .S(_05186_),
    .X(_01149_));
 or4_1 _20299_ (.A(net1302),
    .B(\digitop_pav2.crc_inst.pie_data_en_ff ),
    .C(\digitop_pav2.crc_eval ),
    .D(\digitop_pav2.crc_inst.mctrl_data_en_ff ),
    .X(_05187_));
 and2_1 _20300_ (.A(net1438),
    .B(net1221),
    .X(_00277_));
 nand2_1 _20301_ (.A(net532),
    .B(_11022_),
    .Y(_05188_));
 or3b_1 _20302_ (.A(_05188_),
    .B(net189),
    .C_N(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[0] ),
    .X(_05189_));
 or3b_1 _20303_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[0] ),
    .B(net530),
    .C_N(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[2] ),
    .X(_05190_));
 nor2_1 _20304_ (.A(_11057_),
    .B(_11063_),
    .Y(_05191_));
 or3_1 _20305_ (.A(_11054_),
    .B(_11061_),
    .C(_05191_),
    .X(_05192_));
 a31o_1 _20306_ (.A1(_05189_),
    .A2(_05190_),
    .A3(_05192_),
    .B1(_11042_),
    .X(_05193_));
 or4_1 _20307_ (.A(net532),
    .B(_11022_),
    .C(_11025_),
    .D(_11045_),
    .X(_05194_));
 a21o_1 _20308_ (.A1(_11025_),
    .A2(_11060_),
    .B1(_11061_),
    .X(_05195_));
 and3_1 _20309_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.n_data_valid ),
    .B(_05194_),
    .C(_05195_),
    .X(_05196_));
 o31a_1 _20310_ (.A1(net532),
    .A2(_11039_),
    .A3(_11045_),
    .B1(_11055_),
    .X(_05197_));
 o211ai_4 _20311_ (.A1(_05191_),
    .A2(_05197_),
    .B1(_05196_),
    .C1(_05193_),
    .Y(_05198_));
 inv_2 _20312_ (.A(_05198_),
    .Y(_05199_));
 nor2_1 _20313_ (.A(_11026_),
    .B(_11043_),
    .Y(_05200_));
 a211o_1 _20314_ (.A1(_11048_),
    .A2(_11059_),
    .B1(_05198_),
    .C1(_05200_),
    .X(_05201_));
 nor3_1 _20315_ (.A(net189),
    .B(net191),
    .C(net190),
    .Y(_05202_));
 and2b_1 _20316_ (.A_N(_11042_),
    .B(_05202_),
    .X(_05203_));
 and3b_1 _20317_ (.A_N(net190),
    .B(net191),
    .C(net189),
    .X(_05204_));
 and3_1 _20318_ (.A(net189),
    .B(net191),
    .C(net190),
    .X(_05205_));
 a31o_1 _20319_ (.A1(_11057_),
    .A2(_11061_),
    .A3(_05188_),
    .B1(_05205_),
    .X(_05206_));
 a31o_1 _20320_ (.A1(net529),
    .A2(_11045_),
    .A3(_11063_),
    .B1(_05206_),
    .X(_05207_));
 a21o_1 _20321_ (.A1(_11042_),
    .A2(_05204_),
    .B1(_05207_),
    .X(_05208_));
 o32a_1 _20322_ (.A1(_05201_),
    .A2(_05203_),
    .A3(_05208_),
    .B1(_05199_),
    .B2(net191),
    .X(_01166_));
 a21o_1 _20323_ (.A1(_11042_),
    .A2(_05205_),
    .B1(_05198_),
    .X(_05209_));
 or3b_1 _20324_ (.A(net189),
    .B(net191),
    .C_N(net190),
    .X(_05210_));
 a21oi_1 _20325_ (.A1(net529),
    .A2(_11063_),
    .B1(_05205_),
    .Y(_05211_));
 nor2_1 _20326_ (.A(_11057_),
    .B(_11059_),
    .Y(_05212_));
 mux2_1 _20327_ (.A0(_11025_),
    .A1(_05212_),
    .S(net532),
    .X(_05213_));
 nor2_1 _20328_ (.A(_05202_),
    .B(_05204_),
    .Y(_05214_));
 mux2_1 _20329_ (.A0(_05210_),
    .A1(_05214_),
    .S(_11042_),
    .X(_05215_));
 and3_1 _20330_ (.A(_05211_),
    .B(_05213_),
    .C(_05215_),
    .X(_05216_));
 a2bb2o_1 _20331_ (.A1_N(_05216_),
    .A2_N(_05209_),
    .B1(_05198_),
    .B2(net190),
    .X(_01167_));
 o211a_1 _20332_ (.A1(net532),
    .A2(_11045_),
    .B1(_11057_),
    .C1(_05188_),
    .X(_05217_));
 a311o_1 _20333_ (.A1(net529),
    .A2(_11046_),
    .A3(_11063_),
    .B1(_05204_),
    .C1(_05217_),
    .X(_05218_));
 o21bai_1 _20334_ (.A1(_11042_),
    .A2(_05210_),
    .B1_N(_05218_),
    .Y(_05219_));
 a2bb2o_1 _20335_ (.A1_N(_11043_),
    .A2_N(_11060_),
    .B1(_11048_),
    .B2(_11027_),
    .X(_05220_));
 o32a_1 _20336_ (.A1(_05209_),
    .A2(_05219_),
    .A3(_05220_),
    .B1(_05199_),
    .B2(net189),
    .X(_01168_));
 and2_1 _20337_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[1] ),
    .B(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[0] ),
    .X(_05221_));
 a31oi_1 _20338_ (.A1(_09537_),
    .A2(_11051_),
    .A3(_05221_),
    .B1(_11050_),
    .Y(_05222_));
 nor3b_1 _20339_ (.A(_09565_),
    .B(_05222_),
    .C_N(_09548_),
    .Y(_05223_));
 and2_1 _20340_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[0] ),
    .B(_05223_),
    .X(_05224_));
 nor2_1 _20341_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[0] ),
    .B(_05223_),
    .Y(_05225_));
 nor2_1 _20342_ (.A(_05224_),
    .B(_05225_),
    .Y(_01169_));
 nand2_1 _20343_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[1] ),
    .B(_05224_),
    .Y(_05226_));
 or2_1 _20344_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[1] ),
    .B(_05224_),
    .X(_05227_));
 and2_1 _20345_ (.A(_05226_),
    .B(_05227_),
    .X(_01170_));
 nand2_1 _20346_ (.A(_09563_),
    .B(_05223_),
    .Y(_05228_));
 xnor2_1 _20347_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[2] ),
    .B(_05226_),
    .Y(_01171_));
 or2_1 _20348_ (.A(_07124_),
    .B(_05228_),
    .X(_05229_));
 xnor2_1 _20349_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[3] ),
    .B(_05228_),
    .Y(_01172_));
 xnor2_1 _20350_ (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[4] ),
    .B(_05229_),
    .Y(_01173_));
 mux2_1 _20351_ (.A0(_11050_),
    .A1(net530),
    .S(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[0] ),
    .X(_05230_));
 inv_2 _20352_ (.A(_05230_),
    .Y(_01174_));
 nor2_1 _20353_ (.A(_11050_),
    .B(_05221_),
    .Y(_05231_));
 a22o_1 _20354_ (.A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[1] ),
    .A2(net532),
    .B1(_11044_),
    .B2(_05231_),
    .X(_01175_));
 o21a_1 _20355_ (.A1(net532),
    .A2(_05231_),
    .B1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[2] ),
    .X(_05232_));
 a31o_1 _20356_ (.A1(_07125_),
    .A2(_05221_),
    .A3(_05222_),
    .B1(_05232_),
    .X(_01176_));
 mux2_1 _20357_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[0] ),
    .A1(_11041_),
    .S(net530),
    .X(_01177_));
 mux2_1 _20358_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[0] ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[1] ),
    .S(net531),
    .X(_01178_));
 mux2_1 _20359_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[2] ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[1] ),
    .S(net529),
    .X(_01179_));
 mux2_1 _20360_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[2] ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[3] ),
    .S(net531),
    .X(_01180_));
 mux2_1 _20361_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[3] ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[4] ),
    .S(net531),
    .X(_01181_));
 mux2_1 _20362_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[4] ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[5] ),
    .S(net531),
    .X(_01182_));
 mux2_1 _20363_ (.A0(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[6] ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[5] ),
    .S(net529),
    .X(_01183_));
 o31ai_2 _20364_ (.A1(_08483_),
    .A2(_08520_),
    .A3(net1221),
    .B1(net1439),
    .Y(_05233_));
 mux2_1 _20365_ (.A0(_08519_),
    .A1(\digitop_pav2.crc_inst.mctrl_data_end_ff ),
    .S(_05233_),
    .X(_01184_));
 mux2_1 _20366_ (.A0(\digitop_pav2.crc_eval ),
    .A1(\digitop_pav2.crc_inst.mctrl_data_en_ff ),
    .S(_05233_),
    .X(_01195_));
 nand2_1 _20367_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[1] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[0] ),
    .Y(_05234_));
 nand3_1 _20368_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[1] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[2] ),
    .C(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[0] ),
    .Y(_05235_));
 and2_1 _20369_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[4] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[3] ),
    .X(_05236_));
 and4_1 _20370_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[3] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[1] ),
    .C(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[2] ),
    .D(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[0] ),
    .X(_05237_));
 inv_2 _20371_ (.A(_05237_),
    .Y(_05238_));
 nand2_1 _20372_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[4] ),
    .B(_05237_),
    .Y(_05239_));
 and3_1 _20373_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[5] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[4] ),
    .C(_05237_),
    .X(_05240_));
 inv_2 _20374_ (.A(_05240_),
    .Y(_05241_));
 and2_1 _20375_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[6] ),
    .B(_05240_),
    .X(_05242_));
 inv_2 _20376_ (.A(_05242_),
    .Y(_05243_));
 nand2_1 _20377_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[7] ),
    .B(_05242_),
    .Y(_05244_));
 and3_1 _20378_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[8] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[7] ),
    .C(_05242_),
    .X(_05245_));
 inv_2 _20379_ (.A(_05245_),
    .Y(_05246_));
 nand2_1 _20380_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[0] ),
    .B(net1311),
    .Y(_05247_));
 a21o_1 _20381_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[9] ),
    .A2(_05245_),
    .B1(_05247_),
    .X(_01196_));
 and3_2 _20382_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[9] ),
    .B(net1311),
    .C(_05245_),
    .X(_05248_));
 or2_1 _20383_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[1] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[0] ),
    .X(_05249_));
 a31o_1 _20384_ (.A1(net1311),
    .A2(_05234_),
    .A3(_05249_),
    .B1(_05248_),
    .X(_01197_));
 a21o_1 _20385_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[1] ),
    .A2(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[0] ),
    .B1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[2] ),
    .X(_05250_));
 a31o_1 _20386_ (.A1(net1311),
    .A2(_05235_),
    .A3(_05250_),
    .B1(_05248_),
    .X(_01198_));
 a31o_1 _20387_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[1] ),
    .A2(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[2] ),
    .A3(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[0] ),
    .B1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[3] ),
    .X(_05251_));
 a31o_1 _20388_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.en_pctr ),
    .A2(_05238_),
    .A3(_05251_),
    .B1(_05248_),
    .X(_01199_));
 or2_1 _20389_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[4] ),
    .B(_05237_),
    .X(_05252_));
 a31o_1 _20390_ (.A1(net1311),
    .A2(_05239_),
    .A3(_05252_),
    .B1(_05248_),
    .X(_01200_));
 a21o_1 _20391_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[4] ),
    .A2(_05237_),
    .B1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[5] ),
    .X(_05253_));
 a31o_1 _20392_ (.A1(net1311),
    .A2(_05241_),
    .A3(_05253_),
    .B1(_05248_),
    .X(_01201_));
 or2_1 _20393_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[6] ),
    .B(_05240_),
    .X(_05254_));
 a31o_1 _20394_ (.A1(net1311),
    .A2(_05243_),
    .A3(_05254_),
    .B1(_05248_),
    .X(_01202_));
 or2_1 _20395_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[7] ),
    .B(_05242_),
    .X(_05255_));
 a31o_1 _20396_ (.A1(net1311),
    .A2(_05244_),
    .A3(_05255_),
    .B1(_05248_),
    .X(_01203_));
 a31o_1 _20397_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[7] ),
    .A2(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[6] ),
    .A3(_05240_),
    .B1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[8] ),
    .X(_05256_));
 o211a_1 _20398_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[9] ),
    .A2(_05246_),
    .B1(_05256_),
    .C1(net1311),
    .X(_01204_));
 o21a_1 _20399_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[9] ),
    .A2(_05245_),
    .B1(net1311),
    .X(_01205_));
 mux2_1 _20400_ (.A0(_08487_),
    .A1(\digitop_pav2.crc_inst.dt_tx_en_aux ),
    .S(_05233_),
    .X(_01206_));
 a211o_1 _20401_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[1] ),
    .A2(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[2] ),
    .B1(net1310),
    .C1(_07056_),
    .X(_05257_));
 o211a_1 _20402_ (.A1(_07115_),
    .A2(_05257_),
    .B1(_11105_),
    .C1(_07847_),
    .X(_05258_));
 nand2_1 _20403_ (.A(_07056_),
    .B(_11067_),
    .Y(_05259_));
 a21oi_1 _20404_ (.A1(net1826),
    .A2(_05258_),
    .B1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.en_pctr ),
    .Y(_05260_));
 a21oi_1 _20405_ (.A1(_05258_),
    .A2(_05259_),
    .B1(_05260_),
    .Y(_01207_));
 and3_1 _20406_ (.A(net1326),
    .B(net1325),
    .C(_07855_),
    .X(_05261_));
 nand3_2 _20407_ (.A(net1326),
    .B(net1325),
    .C(_07855_),
    .Y(_05262_));
 nor2_1 _20408_ (.A(net1320),
    .B(_05261_),
    .Y(_05263_));
 nand2_2 _20409_ (.A(_10719_),
    .B(_05262_),
    .Y(_05264_));
 xor2_1 _20410_ (.A(net1108),
    .B(net1096),
    .X(_05265_));
 xnor2_1 _20411_ (.A(net1094),
    .B(_05265_),
    .Y(_05266_));
 xnor2_2 _20412_ (.A(net1134),
    .B(net1121),
    .Y(_05267_));
 xor2_1 _20413_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[0] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[4] ),
    .X(_05268_));
 xor2_2 _20414_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[11] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[12] ),
    .X(_05269_));
 xnor2_1 _20415_ (.A(_05268_),
    .B(_05269_),
    .Y(_05270_));
 xnor2_2 _20416_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[8] ),
    .B(_05269_),
    .Y(_05271_));
 xnor2_1 _20417_ (.A(_05268_),
    .B(_05271_),
    .Y(_05272_));
 xnor2_1 _20418_ (.A(_05266_),
    .B(_05267_),
    .Y(_05273_));
 xnor2_1 _20419_ (.A(_05272_),
    .B(_05273_),
    .Y(_05274_));
 nand2_1 _20420_ (.A(net1107),
    .B(net810),
    .Y(_05275_));
 o22a_1 _20421_ (.A1(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[0] ),
    .A2(net1321),
    .B1(_05264_),
    .B2(_05274_),
    .X(_01208_));
 nand2_1 _20422_ (.A(net1035),
    .B(net809),
    .Y(_05276_));
 nand2_1 _20423_ (.A(net1090),
    .B(net810),
    .Y(_05277_));
 a22o_1 _20424_ (.A1(_07081_),
    .A2(net1090),
    .B1(_05276_),
    .B2(_05277_),
    .X(_05278_));
 xor2_2 _20425_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[13] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[9] ),
    .X(_05279_));
 xnor2_1 _20426_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[12] ),
    .B(_05279_),
    .Y(_05280_));
 xor2_2 _20427_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[1] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[5] ),
    .X(_05281_));
 xnor2_1 _20428_ (.A(net1131),
    .B(_05281_),
    .Y(_05282_));
 xnor2_1 _20429_ (.A(_05280_),
    .B(_05282_),
    .Y(_05283_));
 xor2_1 _20430_ (.A(net1118),
    .B(net1103),
    .X(_05284_));
 nand2_1 _20431_ (.A(net1104),
    .B(net809),
    .Y(_05285_));
 nand2_1 _20432_ (.A(net810),
    .B(_05284_),
    .Y(_05286_));
 xnor2_1 _20433_ (.A(_05283_),
    .B(_05286_),
    .Y(_05287_));
 xnor2_1 _20434_ (.A(_05278_),
    .B(_05287_),
    .Y(_05288_));
 a22o_1 _20435_ (.A1(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[1] ),
    .A2(net1320),
    .B1(_05263_),
    .B2(_05288_),
    .X(_01209_));
 xnor2_1 _20436_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[13] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[14] ),
    .Y(_05289_));
 xnor2_1 _20437_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[10] ),
    .B(_05289_),
    .Y(_05290_));
 xor2_2 _20438_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[2] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[6] ),
    .X(_05291_));
 xnor2_1 _20439_ (.A(_05290_),
    .B(_05291_),
    .Y(_05292_));
 xor2_2 _20440_ (.A(net1091),
    .B(net1087),
    .X(_05293_));
 xnor2_4 _20441_ (.A(net1099),
    .B(_05293_),
    .Y(_05294_));
 xor2_2 _20442_ (.A(net1128),
    .B(net1115),
    .X(_05295_));
 xnor2_1 _20443_ (.A(_05294_),
    .B(_05295_),
    .Y(_05296_));
 and2_1 _20444_ (.A(_05292_),
    .B(_05296_),
    .X(_05297_));
 nor2_1 _20445_ (.A(_05292_),
    .B(_05296_),
    .Y(_05298_));
 nand2_1 _20446_ (.A(net809),
    .B(_05295_),
    .Y(_05299_));
 o32a_1 _20447_ (.A1(_05264_),
    .A2(_05297_),
    .A3(_05298_),
    .B1(net1321),
    .B2(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[2] ),
    .X(_01210_));
 nand2_1 _20448_ (.A(net1111),
    .B(net809),
    .Y(_05300_));
 xor2_2 _20449_ (.A(net1083),
    .B(net1087),
    .X(_05301_));
 xnor2_1 _20450_ (.A(net1096),
    .B(_05301_),
    .Y(_05302_));
 nand2_1 _20451_ (.A(net809),
    .B(_05302_),
    .Y(_05303_));
 o22a_1 _20452_ (.A1(_05300_),
    .A2(_05302_),
    .B1(_05303_),
    .B2(net1111),
    .X(_05304_));
 nand2_1 _20453_ (.A(net1124),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[15] ),
    .Y(_05305_));
 or2_1 _20454_ (.A(net1124),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[15] ),
    .X(_05306_));
 xor2_1 _20455_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[3] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[7] ),
    .X(_05307_));
 xnor2_1 _20456_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[11] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[14] ),
    .Y(_05308_));
 xnor2_1 _20457_ (.A(_05307_),
    .B(_05308_),
    .Y(_05309_));
 a21oi_1 _20458_ (.A1(_05305_),
    .A2(_05306_),
    .B1(_05309_),
    .Y(_05310_));
 a31o_1 _20459_ (.A1(_05305_),
    .A2(_05306_),
    .A3(_05309_),
    .B1(_05310_),
    .X(_05311_));
 xnor2_1 _20460_ (.A(_05304_),
    .B(_05311_),
    .Y(_05312_));
 a22o_1 _20461_ (.A1(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[3] ),
    .A2(net1320),
    .B1(_05263_),
    .B2(_05312_),
    .X(_01211_));
 nand2_1 _20462_ (.A(net1084),
    .B(net1095),
    .Y(_05313_));
 or2_1 _20463_ (.A(net1083),
    .B(net1094),
    .X(_05314_));
 nand2_1 _20464_ (.A(_05313_),
    .B(_05314_),
    .Y(_05315_));
 nand2_1 _20465_ (.A(net810),
    .B(_05315_),
    .Y(_05316_));
 o22a_1 _20466_ (.A1(_05275_),
    .A2(_05315_),
    .B1(_05316_),
    .B2(net1108),
    .X(_05317_));
 nand2_1 _20467_ (.A(net1121),
    .B(net810),
    .Y(_05318_));
 xor2_1 _20468_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[4] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[8] ),
    .X(_05319_));
 xor2_1 _20469_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[12] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[15] ),
    .X(_05320_));
 xnor2_1 _20470_ (.A(_05319_),
    .B(_05320_),
    .Y(_05321_));
 xnor2_1 _20471_ (.A(_05318_),
    .B(_05321_),
    .Y(_05322_));
 xnor2_1 _20472_ (.A(_05317_),
    .B(_05322_),
    .Y(_05323_));
 o22a_1 _20473_ (.A1(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[4] ),
    .A2(net1321),
    .B1(_05264_),
    .B2(_05323_),
    .X(_01212_));
 xnor2_1 _20474_ (.A(net1096),
    .B(_05284_),
    .Y(_05324_));
 nand2_1 _20475_ (.A(net810),
    .B(_05324_),
    .Y(_05325_));
 xnor2_1 _20476_ (.A(_05278_),
    .B(_05325_),
    .Y(_05326_));
 xor2_1 _20477_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[8] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[5] ),
    .X(_05327_));
 xnor2_1 _20478_ (.A(_05279_),
    .B(_05327_),
    .Y(_05328_));
 xnor2_1 _20479_ (.A(_05270_),
    .B(_05328_),
    .Y(_05329_));
 nor2_1 _20480_ (.A(net1320),
    .B(net809),
    .Y(_05330_));
 a211oi_1 _20481_ (.A1(net1134),
    .A2(net810),
    .B1(_05329_),
    .C1(_05330_),
    .Y(_05331_));
 a31o_1 _20482_ (.A1(net1134),
    .A2(net810),
    .A3(_05329_),
    .B1(_05331_),
    .X(_05332_));
 xor2_1 _20483_ (.A(net1121),
    .B(net1108),
    .X(_05333_));
 nand2_1 _20484_ (.A(net810),
    .B(_05333_),
    .Y(_05334_));
 xnor2_1 _20485_ (.A(_05332_),
    .B(_05334_),
    .Y(_05335_));
 xnor2_1 _20486_ (.A(_05326_),
    .B(_05335_),
    .Y(_05336_));
 mux2_1 _20487_ (.A0(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[5] ),
    .A1(_05336_),
    .S(net1321),
    .X(_01213_));
 xnor2_1 _20488_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[10] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[9] ),
    .Y(_05337_));
 xnor2_1 _20489_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[10] ),
    .B(_05279_),
    .Y(_05338_));
 xor2_1 _20490_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[12] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[6] ),
    .X(_05339_));
 xnor2_1 _20491_ (.A(_05281_),
    .B(_05339_),
    .Y(_05340_));
 xor2_2 _20492_ (.A(net1131),
    .B(net1118),
    .X(_05341_));
 xnor2_1 _20493_ (.A(net1094),
    .B(_05341_),
    .Y(_05342_));
 xnor2_1 _20494_ (.A(net1115),
    .B(net1104),
    .Y(_05343_));
 xnor2_1 _20495_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[14] ),
    .B(_05343_),
    .Y(_05344_));
 xnor2_1 _20496_ (.A(_05338_),
    .B(_05340_),
    .Y(_05345_));
 xnor2_1 _20497_ (.A(_05294_),
    .B(_05342_),
    .Y(_05346_));
 xnor2_1 _20498_ (.A(_05345_),
    .B(_05346_),
    .Y(_05347_));
 xnor2_1 _20499_ (.A(_05344_),
    .B(_05347_),
    .Y(_05348_));
 o22a_1 _20500_ (.A1(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[6] ),
    .A2(net1321),
    .B1(_05264_),
    .B2(_05348_),
    .X(_01214_));
 xor2_1 _20501_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[14] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[15] ),
    .X(_05349_));
 xor2_1 _20502_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[11] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[13] ),
    .X(_05350_));
 xnor2_1 _20503_ (.A(_05349_),
    .B(_05350_),
    .Y(_05351_));
 xor2_1 _20504_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[10] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[7] ),
    .X(_05352_));
 xor2_1 _20505_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[10] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[6] ),
    .X(_05353_));
 xnor2_1 _20506_ (.A(_05291_),
    .B(_05352_),
    .Y(_05354_));
 xnor2_1 _20507_ (.A(_05351_),
    .B(_05354_),
    .Y(_05355_));
 nor2_1 _20508_ (.A(_05330_),
    .B(_05355_),
    .Y(_05356_));
 mux2_1 _20509_ (.A0(_05355_),
    .A1(_05356_),
    .S(_05299_),
    .X(_05357_));
 nand2_1 _20510_ (.A(net1100),
    .B(_05262_),
    .Y(_05358_));
 o22a_1 _20511_ (.A1(net1100),
    .A2(_05303_),
    .B1(_05358_),
    .B2(_05302_),
    .X(_05359_));
 a22o_1 _20512_ (.A1(net1111),
    .A2(net1091),
    .B1(_05277_),
    .B2(_05300_),
    .X(_05360_));
 xnor2_1 _20513_ (.A(_05359_),
    .B(_05360_),
    .Y(_05361_));
 nor2_1 _20514_ (.A(_05357_),
    .B(_05361_),
    .Y(_05362_));
 a21o_1 _20515_ (.A1(_05357_),
    .A2(_05361_),
    .B1(net1320),
    .X(_05363_));
 a2bb2o_1 _20516_ (.A1_N(_05362_),
    .A2_N(_05363_),
    .B1(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[7] ),
    .B2(net1320),
    .X(_01215_));
 nand2_1 _20517_ (.A(net1124),
    .B(net809),
    .Y(_05364_));
 xnor2_1 _20518_ (.A(_05307_),
    .B(_05349_),
    .Y(_05365_));
 xnor2_1 _20519_ (.A(_05271_),
    .B(_05365_),
    .Y(_05366_));
 o21ai_1 _20520_ (.A1(net1320),
    .A2(net809),
    .B1(_05366_),
    .Y(_05367_));
 mux2_1 _20521_ (.A0(_05366_),
    .A1(_05367_),
    .S(_05364_),
    .X(_05368_));
 o22a_1 _20522_ (.A1(_05276_),
    .A2(_05302_),
    .B1(_05303_),
    .B2(net1035),
    .X(_05369_));
 a22o_1 _20523_ (.A1(net1111),
    .A2(net1108),
    .B1(_05275_),
    .B2(_05300_),
    .X(_05370_));
 xnor2_1 _20524_ (.A(_05369_),
    .B(_05370_),
    .Y(_05371_));
 nor2_1 _20525_ (.A(_05368_),
    .B(_05371_),
    .Y(_05372_));
 a21o_1 _20526_ (.A1(_05368_),
    .A2(_05371_),
    .B1(_10720_),
    .X(_05373_));
 o22a_1 _20527_ (.A1(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[8] ),
    .A2(net1321),
    .B1(_05372_),
    .B2(_05373_),
    .X(_01216_));
 o22a_1 _20528_ (.A1(_05277_),
    .A2(_05315_),
    .B1(_05316_),
    .B2(net1090),
    .X(_05374_));
 xnor2_1 _20529_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[15] ),
    .B(_05319_),
    .Y(_05375_));
 xnor2_1 _20530_ (.A(_05280_),
    .B(_05375_),
    .Y(_05376_));
 xnor2_1 _20531_ (.A(_05374_),
    .B(_05376_),
    .Y(_05377_));
 xnor2_1 _20532_ (.A(_05285_),
    .B(_05334_),
    .Y(_05378_));
 nor2_1 _20533_ (.A(_05377_),
    .B(_05378_),
    .Y(_05379_));
 a21o_1 _20534_ (.A1(_05377_),
    .A2(_05378_),
    .B1(_05264_),
    .X(_05380_));
 o22a_1 _20535_ (.A1(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[9] ),
    .A2(net1321),
    .B1(_05379_),
    .B2(_05380_),
    .X(_01217_));
 xor2_1 _20536_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[5] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[14] ),
    .X(_05381_));
 xnor2_1 _20537_ (.A(_05338_),
    .B(_05381_),
    .Y(_05382_));
 o22ai_1 _20538_ (.A1(_05261_),
    .A2(_05294_),
    .B1(_05330_),
    .B2(_05382_),
    .Y(_05383_));
 o31ai_1 _20539_ (.A1(_05261_),
    .A2(_05294_),
    .A3(_05382_),
    .B1(_05383_),
    .Y(_05384_));
 xnor2_1 _20540_ (.A(_05286_),
    .B(_05384_),
    .Y(_05385_));
 mux2_1 _20541_ (.A0(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[10] ),
    .A1(_05385_),
    .S(net1321),
    .X(_01218_));
 xor2_1 _20542_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[10] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[11] ),
    .X(_05386_));
 xnor2_1 _20543_ (.A(_05308_),
    .B(_05353_),
    .Y(_05387_));
 nand2_1 _20544_ (.A(net1115),
    .B(net809),
    .Y(_05388_));
 xnor2_1 _20545_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[15] ),
    .B(_05388_),
    .Y(_05389_));
 xnor2_1 _20546_ (.A(_05359_),
    .B(_05389_),
    .Y(_05390_));
 xnor2_1 _20547_ (.A(_05387_),
    .B(_05390_),
    .Y(_05391_));
 a22o_1 _20548_ (.A1(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[11] ),
    .A2(net1320),
    .B1(_05263_),
    .B2(_05391_),
    .X(_01219_));
 xor2_1 _20549_ (.A(net1134),
    .B(net1111),
    .X(_05392_));
 xnor2_1 _20550_ (.A(net1084),
    .B(_05333_),
    .Y(_05393_));
 xnor2_1 _20551_ (.A(_05392_),
    .B(_05393_),
    .Y(_05394_));
 xnor2_1 _20552_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[7] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[0] ),
    .Y(_05395_));
 xnor2_1 _20553_ (.A(_05375_),
    .B(_05395_),
    .Y(_05396_));
 nor2_1 _20554_ (.A(_05394_),
    .B(_05396_),
    .Y(_05397_));
 and2_1 _20555_ (.A(_05394_),
    .B(_05396_),
    .X(_05398_));
 o32a_1 _20556_ (.A1(_05264_),
    .A2(_05397_),
    .A3(_05398_),
    .B1(net1321),
    .B2(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[12] ),
    .X(_01220_));
 nand2_1 _20557_ (.A(net810),
    .B(_05341_),
    .Y(_05399_));
 xor2_1 _20558_ (.A(_05281_),
    .B(_05399_),
    .X(_05400_));
 a22o_1 _20559_ (.A1(net1108),
    .A2(net1104),
    .B1(_05275_),
    .B2(_05285_),
    .X(_05401_));
 xnor2_1 _20560_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[8] ),
    .B(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[9] ),
    .Y(_05402_));
 xnor2_1 _20561_ (.A(_05401_),
    .B(_05402_),
    .Y(_05403_));
 or2_1 _20562_ (.A(_05400_),
    .B(_05403_),
    .X(_05404_));
 nand2_1 _20563_ (.A(_05400_),
    .B(_05403_),
    .Y(_05405_));
 a32o_1 _20564_ (.A1(_05263_),
    .A2(_05404_),
    .A3(_05405_),
    .B1(net1320),
    .B2(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[13] ),
    .X(_01221_));
 a22o_1 _20565_ (.A1(net1104),
    .A2(net1099),
    .B1(_05285_),
    .B2(_05358_),
    .X(_05406_));
 xnor2_1 _20566_ (.A(_05291_),
    .B(_05337_),
    .Y(_05407_));
 xnor2_1 _20567_ (.A(_05299_),
    .B(_05407_),
    .Y(_05408_));
 xnor2_1 _20568_ (.A(_05406_),
    .B(_05408_),
    .Y(_05409_));
 a22o_1 _20569_ (.A1(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[14] ),
    .A2(net1320),
    .B1(_05263_),
    .B2(_05409_),
    .X(_01222_));
 nand2_1 _20570_ (.A(_07080_),
    .B(net809),
    .Y(_05410_));
 mux2_1 _20571_ (.A0(_05410_),
    .A1(_05358_),
    .S(net1096),
    .X(_05411_));
 xor2_1 _20572_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[7] ),
    .B(_05300_),
    .X(_05412_));
 xnor2_1 _20573_ (.A(_05411_),
    .B(_05412_),
    .Y(_05413_));
 xnor2_1 _20574_ (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[3] ),
    .B(_05386_),
    .Y(_05414_));
 xnor2_1 _20575_ (.A(_05364_),
    .B(_05414_),
    .Y(_05415_));
 xnor2_1 _20576_ (.A(_05413_),
    .B(_05415_),
    .Y(_05416_));
 o22a_1 _20577_ (.A1(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[15] ),
    .A2(_10719_),
    .B1(_05264_),
    .B2(_05416_),
    .X(_01223_));
 or2_1 _20578_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[1] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[2] ),
    .X(_05417_));
 or3_1 _20579_ (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[5] ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[6] ),
    .C(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[9] ),
    .X(_05418_));
 a2111oi_1 _20580_ (.A1(_05236_),
    .A2(_05417_),
    .B1(_05418_),
    .C1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[7] ),
    .D1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[8] ),
    .Y(_05419_));
 a21boi_1 _20581_ (.A1(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[0] ),
    .A2(_05236_),
    .B1_N(_05419_),
    .Y(_05420_));
 and2_1 _20582_ (.A(\digitop_pav2.cal_inst.calx_mux.dtest_trim_0_i ),
    .B(_05420_),
    .X(_05421_));
 and2b_1 _20583_ (.A_N(_05421_),
    .B(net1306),
    .X(_05422_));
 or2_1 _20584_ (.A(net1826),
    .B(_05257_),
    .X(_05423_));
 nor2_1 _20585_ (.A(net1826),
    .B(_05257_),
    .Y(_05424_));
 a31o_1 _20586_ (.A1(\digitop_pav2.cal_inst.calx_mux.dtest_trim_2_i ),
    .A2(\digitop_pav2.cal_inst.calx_mux.dtest_trim_1_i ),
    .A3(\digitop_pav2.cal_inst.calx_mux.dtest_trim_0_i ),
    .B1(_05423_),
    .X(_05425_));
 o21a_1 _20587_ (.A1(net1306),
    .A2(_05423_),
    .B1(_05425_),
    .X(_05426_));
 o22a_1 _20588_ (.A1(\digitop_pav2.cal_inst.calx_mux.dtest_trim_0_i ),
    .A2(_05420_),
    .B1(_05422_),
    .B2(_05426_),
    .X(_05427_));
 nor2_1 _20589_ (.A(\digitop_pav2.cal_inst.calx_mux.dtest_trim_0_i ),
    .B(net1306),
    .Y(_05428_));
 o21a_1 _20590_ (.A1(\digitop_pav2.cal_inst.calx_mux.dtest_trim_2_i ),
    .A2(\digitop_pav2.cal_inst.calx_mux.dtest_trim_1_i ),
    .B1(_05428_),
    .X(_05429_));
 o22a_1 _20591_ (.A1(\digitop_pav2.cal_inst.calx_mux.dtest_trim_0_i ),
    .A2(_05424_),
    .B1(_05427_),
    .B2(_05429_),
    .X(_01224_));
 o221a_1 _20592_ (.A1(\digitop_pav2.cal_inst.calx_mux.dtest_trim_2_i ),
    .A2(\digitop_pav2.cal_inst.calx_mux.dtest_trim_0_i ),
    .B1(_05421_),
    .B2(_05428_),
    .C1(_07116_),
    .X(_05430_));
 a2bb2o_1 _20593_ (.A1_N(_05425_),
    .A2_N(_05430_),
    .B1(_07116_),
    .B2(_05423_),
    .X(_05431_));
 o31ai_1 _20594_ (.A1(_07116_),
    .A2(_05421_),
    .A3(_05428_),
    .B1(_05431_),
    .Y(_01225_));
 a21oi_1 _20595_ (.A1(\digitop_pav2.cal_inst.calx_mux.dtest_trim_1_i ),
    .A2(_05421_),
    .B1(\digitop_pav2.cal_inst.calx_mux.dtest_trim_2_i ),
    .Y(_05432_));
 a21oi_1 _20596_ (.A1(_07116_),
    .A2(_05428_),
    .B1(_05432_),
    .Y(_05433_));
 o22a_1 _20597_ (.A1(\digitop_pav2.cal_inst.calx_mux.dtest_trim_2_i ),
    .A2(_05424_),
    .B1(_05425_),
    .B2(_05433_),
    .X(_01226_));
 o21a_1 _20598_ (.A1(\digitop_pav2.boot_inst.boot_ctrl0.prev_busy ),
    .A2(net1445),
    .B1(_10718_),
    .X(_01227_));
 a21oi_1 _20599_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[2] ),
    .A2(_10742_),
    .B1(net464),
    .Y(_05434_));
 inv_2 _20600_ (.A(net346),
    .Y(_05435_));
 and2_1 _20601_ (.A(net390),
    .B(_05435_),
    .X(_05436_));
 nand2_1 _20602_ (.A(net390),
    .B(_05435_),
    .Y(_05437_));
 a21o_1 _20603_ (.A1(net455),
    .A2(_07227_),
    .B1(net301),
    .X(_05438_));
 o21ai_1 _20604_ (.A1(_07546_),
    .A2(_02559_),
    .B1(_07108_),
    .Y(_05439_));
 nor2_1 _20605_ (.A(_07548_),
    .B(_03001_),
    .Y(_05440_));
 o2bb2a_1 _20606_ (.A1_N(net1135),
    .A2_N(_05439_),
    .B1(_05440_),
    .B2(_02559_),
    .X(_05441_));
 nor2_2 _20607_ (.A(net455),
    .B(_05441_),
    .Y(_05442_));
 a31o_1 _20608_ (.A1(net455),
    .A2(_07197_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key2_r[0] ),
    .B1(_05442_),
    .X(_05443_));
 a22o_1 _20609_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[0] ),
    .A2(_05438_),
    .B1(_05443_),
    .B2(net303),
    .X(_01228_));
 a21o_1 _20610_ (.A1(net452),
    .A2(_07228_),
    .B1(net302),
    .X(_05444_));
 a22o_1 _20611_ (.A1(net1132),
    .A2(net714),
    .B1(_05440_),
    .B2(net1255),
    .X(_05445_));
 o211a_2 _20612_ (.A1(net1132),
    .A2(_07546_),
    .B1(_05445_),
    .C1(net412),
    .X(_05446_));
 a31o_1 _20613_ (.A1(net452),
    .A2(_07195_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key2_r[1] ),
    .B1(_05446_),
    .X(_05447_));
 a22o_1 _20614_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[1] ),
    .A2(_05444_),
    .B1(_05447_),
    .B2(net304),
    .X(_01229_));
 a21o_1 _20615_ (.A1(net450),
    .A2(_07229_),
    .B1(net302),
    .X(_05448_));
 a21oi_1 _20616_ (.A1(_08118_),
    .A2(_02270_),
    .B1(_07548_),
    .Y(_05449_));
 o2bb2a_2 _20617_ (.A1_N(net1130),
    .A2_N(_05439_),
    .B1(_05449_),
    .B2(_02559_),
    .X(_05450_));
 nor2_2 _20618_ (.A(net451),
    .B(_05450_),
    .Y(_05451_));
 a31o_1 _20619_ (.A1(net450),
    .A2(_07199_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key2_r[2] ),
    .B1(_05451_),
    .X(_05452_));
 a22o_1 _20620_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[2] ),
    .A2(_05448_),
    .B1(_05452_),
    .B2(net304),
    .X(_01230_));
 a21o_1 _20621_ (.A1(net456),
    .A2(_07230_),
    .B1(net302),
    .X(_05453_));
 nor2_2 _20622_ (.A(_07475_),
    .B(_07548_),
    .Y(_05454_));
 a22o_1 _20623_ (.A1(net1126),
    .A2(net714),
    .B1(_05454_),
    .B2(net1255),
    .X(_05455_));
 o211a_2 _20624_ (.A1(net1036),
    .A2(net1126),
    .B1(net412),
    .C1(_05455_),
    .X(_05456_));
 a31o_1 _20625_ (.A1(net456),
    .A2(_07201_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key2_r[3] ),
    .B1(_05456_),
    .X(_05457_));
 a22o_1 _20626_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[3] ),
    .A2(_05453_),
    .B1(_05457_),
    .B2(net304),
    .X(_01231_));
 a21o_1 _20627_ (.A1(net465),
    .A2(_07231_),
    .B1(net302),
    .X(_05458_));
 a31o_2 _20628_ (.A1(net1155),
    .A2(net1255),
    .A3(_05454_),
    .B1(net714),
    .X(_05459_));
 and3_2 _20629_ (.A(net1123),
    .B(net409),
    .C(_05459_),
    .X(_05460_));
 a31o_1 _20630_ (.A1(net465),
    .A2(_07203_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key2_r[4] ),
    .B1(_05460_),
    .X(_05461_));
 a22o_1 _20631_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[4] ),
    .A2(_05458_),
    .B1(_05461_),
    .B2(net304),
    .X(_01232_));
 a21o_1 _20632_ (.A1(net465),
    .A2(_07232_),
    .B1(net302),
    .X(_05462_));
 a31o_1 _20633_ (.A1(net1155),
    .A2(_07077_),
    .A3(_05454_),
    .B1(_02559_),
    .X(_05463_));
 nand2_1 _20634_ (.A(net1120),
    .B(net714),
    .Y(_05464_));
 a21oi_4 _20635_ (.A1(_05463_),
    .A2(_05464_),
    .B1(net458),
    .Y(_05465_));
 a31o_1 _20636_ (.A1(net465),
    .A2(_07205_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key2_r[5] ),
    .B1(_05465_),
    .X(_05466_));
 a22o_1 _20637_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[5] ),
    .A2(_05462_),
    .B1(_05466_),
    .B2(net304),
    .X(_01233_));
 a21o_1 _20638_ (.A1(net451),
    .A2(_07233_),
    .B1(net302),
    .X(_05467_));
 a31o_1 _20639_ (.A1(net1155),
    .A2(_07078_),
    .A3(_05454_),
    .B1(_02559_),
    .X(_05468_));
 nand2_1 _20640_ (.A(net1117),
    .B(net714),
    .Y(_05469_));
 a21oi_4 _20641_ (.A1(_05468_),
    .A2(_05469_),
    .B1(net458),
    .Y(_05470_));
 a31o_1 _20642_ (.A1(net451),
    .A2(_07207_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key2_r[6] ),
    .B1(_05470_),
    .X(_05471_));
 a22o_1 _20643_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[6] ),
    .A2(_05467_),
    .B1(_05471_),
    .B2(net304),
    .X(_01234_));
 a21o_1 _20644_ (.A1(net445),
    .A2(_07234_),
    .B1(net301),
    .X(_05472_));
 and3_2 _20645_ (.A(net1114),
    .B(net407),
    .C(_05459_),
    .X(_05473_));
 a31o_1 _20646_ (.A1(net445),
    .A2(_07209_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key2_r[7] ),
    .B1(_05473_),
    .X(_05474_));
 a22o_1 _20647_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[7] ),
    .A2(_05472_),
    .B1(_05474_),
    .B2(net303),
    .X(_01235_));
 a21o_1 _20648_ (.A1(net447),
    .A2(_07171_),
    .B1(net301),
    .X(_05475_));
 o2bb2a_1 _20649_ (.A1_N(net1110),
    .A2_N(_05459_),
    .B1(_07549_),
    .B2(_07477_),
    .X(_05476_));
 nor2_2 _20650_ (.A(net461),
    .B(_05476_),
    .Y(_05477_));
 a31o_1 _20651_ (.A1(net447),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[8] ),
    .A3(_07172_),
    .B1(_05477_),
    .X(_05478_));
 a22o_1 _20652_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[8] ),
    .A2(_05475_),
    .B1(_05478_),
    .B2(net303),
    .X(_01236_));
 a21o_1 _20653_ (.A1(net443),
    .A2(_07173_),
    .B1(net301),
    .X(_05479_));
 and3_2 _20654_ (.A(net1106),
    .B(net407),
    .C(_05459_),
    .X(_05480_));
 a31o_1 _20655_ (.A1(net443),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[9] ),
    .A3(_07174_),
    .B1(_05480_),
    .X(_05481_));
 a22o_1 _20656_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[9] ),
    .A2(_05479_),
    .B1(_05481_),
    .B2(net303),
    .X(_01237_));
 a21o_1 _20657_ (.A1(net447),
    .A2(_07175_),
    .B1(net301),
    .X(_05482_));
 o2bb2a_1 _20658_ (.A1_N(net1102),
    .A2_N(_05459_),
    .B1(_07549_),
    .B2(_02270_),
    .X(_05483_));
 nor2_2 _20659_ (.A(net447),
    .B(_05483_),
    .Y(_05484_));
 a31o_1 _20660_ (.A1(net447),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[10] ),
    .A3(_07176_),
    .B1(_05484_),
    .X(_05485_));
 a22o_1 _20661_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[10] ),
    .A2(_05482_),
    .B1(_05485_),
    .B2(net303),
    .X(_01238_));
 a21o_1 _20662_ (.A1(net460),
    .A2(_07177_),
    .B1(net301),
    .X(_05486_));
 a21oi_1 _20663_ (.A1(_07025_),
    .A2(net1036),
    .B1(_07548_),
    .Y(_05487_));
 o2bb2a_2 _20664_ (.A1_N(net1098),
    .A2_N(_05439_),
    .B1(_05487_),
    .B2(_02559_),
    .X(_05488_));
 nor2_2 _20665_ (.A(net461),
    .B(_05488_),
    .Y(_05489_));
 a31o_1 _20666_ (.A1(net460),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[11] ),
    .A3(_07178_),
    .B1(_05489_),
    .X(_05490_));
 a22o_1 _20667_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[11] ),
    .A2(_05486_),
    .B1(_05490_),
    .B2(net303),
    .X(_01239_));
 a21o_1 _20668_ (.A1(net460),
    .A2(_07179_),
    .B1(net301),
    .X(_05491_));
 o21a_1 _20669_ (.A1(net1036),
    .A2(net1035),
    .B1(_05454_),
    .X(_05492_));
 o22a_2 _20670_ (.A1(net1035),
    .A2(_07108_),
    .B1(_02559_),
    .B2(_05492_),
    .X(_05493_));
 nor2_2 _20671_ (.A(net461),
    .B(_05493_),
    .Y(_05494_));
 a31o_1 _20672_ (.A1(net460),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[12] ),
    .A3(_07180_),
    .B1(_05494_),
    .X(_05495_));
 a22o_1 _20673_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[12] ),
    .A2(_05491_),
    .B1(_05495_),
    .B2(net303),
    .X(_01240_));
 a21o_1 _20674_ (.A1(net449),
    .A2(_07181_),
    .B1(net301),
    .X(_05496_));
 a31o_1 _20675_ (.A1(net1155),
    .A2(_07082_),
    .A3(_05454_),
    .B1(_02559_),
    .X(_05497_));
 nand2_1 _20676_ (.A(net1093),
    .B(net714),
    .Y(_05498_));
 a21oi_4 _20677_ (.A1(_05497_),
    .A2(_05498_),
    .B1(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[5] ),
    .Y(_05499_));
 a31o_1 _20678_ (.A1(net462),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[13] ),
    .A3(_07182_),
    .B1(_05499_),
    .X(_05500_));
 a22o_1 _20679_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[13] ),
    .A2(_05496_),
    .B1(_05500_),
    .B2(net303),
    .X(_01241_));
 a21o_1 _20680_ (.A1(net442),
    .A2(_07183_),
    .B1(net301),
    .X(_05501_));
 a31o_1 _20681_ (.A1(net1155),
    .A2(_07083_),
    .A3(_05454_),
    .B1(_02559_),
    .X(_05502_));
 nand2_1 _20682_ (.A(net1089),
    .B(net714),
    .Y(_05503_));
 a21oi_4 _20683_ (.A1(_05502_),
    .A2(_05503_),
    .B1(net457),
    .Y(_05504_));
 a31o_1 _20684_ (.A1(net442),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[14] ),
    .A3(_07184_),
    .B1(_05504_),
    .X(_05505_));
 a22o_1 _20685_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[14] ),
    .A2(_05501_),
    .B1(_05505_),
    .B2(net303),
    .X(_01242_));
 a21o_1 _20686_ (.A1(net442),
    .A2(_07185_),
    .B1(net301),
    .X(_05506_));
 and3_2 _20687_ (.A(net1086),
    .B(net407),
    .C(_05459_),
    .X(_05507_));
 a31o_1 _20688_ (.A1(net442),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[15] ),
    .A3(_07186_),
    .B1(_05507_),
    .X(_05508_));
 a22o_1 _20689_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key0_r[15] ),
    .A2(_05506_),
    .B1(_05508_),
    .B2(net303),
    .X(_01243_));
 a21o_1 _20690_ (.A1(_07832_),
    .A2(_10726_),
    .B1(net1326),
    .X(_05509_));
 nand3_1 _20691_ (.A(\digitop_pav2.boot_inst.boot_proc0.proc_stage[0] ),
    .B(_07832_),
    .C(_10726_),
    .Y(_05510_));
 nand2_1 _20692_ (.A(_05509_),
    .B(_05510_),
    .Y(_01244_));
 xnor2_1 _20693_ (.A(\digitop_pav2.boot_inst.boot_proc0.proc_stage[1] ),
    .B(_05509_),
    .Y(_01245_));
 a21o_1 _20694_ (.A1(\digitop_pav2.boot_inst.boot_ctrl0.act_state_i ),
    .A2(net1317),
    .B1(_07835_),
    .X(_01246_));
 mux2_1 _20695_ (.A0(net1132),
    .A1(net1324),
    .S(net1316),
    .X(_01247_));
 mux2_1 _20696_ (.A0(net1130),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[1] ),
    .S(net1316),
    .X(_01248_));
 mux2_1 _20697_ (.A0(net1126),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[2] ),
    .S(net1316),
    .X(_01249_));
 mux2_1 _20698_ (.A0(net1121),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[3] ),
    .S(net1317),
    .X(_01250_));
 mux2_1 _20699_ (.A0(net1118),
    .A1(net1323),
    .S(net1317),
    .X(_01251_));
 mux2_1 _20700_ (.A0(net1117),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[5] ),
    .S(net1316),
    .X(_01252_));
 mux2_1 _20701_ (.A0(net1112),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[6] ),
    .S(net1316),
    .X(_01253_));
 mux2_1 _20702_ (.A0(net1110),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[7] ),
    .S(net1316),
    .X(_01254_));
 mux2_1 _20703_ (.A0(net1103),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[8] ),
    .S(net1317),
    .X(_01255_));
 mux2_1 _20704_ (.A0(net1102),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[9] ),
    .S(net1316),
    .X(_01256_));
 mux2_1 _20705_ (.A0(net1098),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[10] ),
    .S(net1316),
    .X(_01257_));
 mux2_1 _20706_ (.A0(net1094),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[11] ),
    .S(net1316),
    .X(_01258_));
 mux2_1 _20707_ (.A0(net1090),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_fg[12] ),
    .S(net1317),
    .X(_01259_));
 mux2_1 _20708_ (.A0(net1087),
    .A1(\digitop_pav2.access_inst.access_check0.fg_i[13] ),
    .S(net1316),
    .X(_01260_));
 and2_1 _20709_ (.A(net1322),
    .B(_07826_),
    .X(_05511_));
 nor2_1 _20710_ (.A(_07082_),
    .B(_07832_),
    .Y(_05512_));
 or4b_1 _20711_ (.A(net1326),
    .B(net1091),
    .C(net1087),
    .D_N(\digitop_pav2.boot_inst.boot_proc0.proc_stage[1] ),
    .X(_05513_));
 or2_1 _20712_ (.A(_05313_),
    .B(_05513_),
    .X(_05514_));
 and4_1 _20713_ (.A(net1325),
    .B(net1083),
    .C(net1112),
    .D(net1104),
    .X(_05515_));
 nand2_1 _20714_ (.A(net1134),
    .B(_05515_),
    .Y(_05516_));
 or4_1 _20715_ (.A(net1325),
    .B(net1083),
    .C(net1111),
    .D(net1104),
    .X(_05517_));
 o21a_1 _20716_ (.A1(net1134),
    .A2(_05517_),
    .B1(_07082_),
    .X(_05518_));
 or4_1 _20717_ (.A(net1131),
    .B(net1124),
    .C(net1121),
    .D(net1118),
    .X(_05519_));
 or4b_1 _20718_ (.A(net1128),
    .B(net1115),
    .C(net1108),
    .D_N(net1326),
    .X(_05520_));
 or4_1 _20719_ (.A(net1100),
    .B(net1094),
    .C(_07083_),
    .D(_05520_),
    .X(_05521_));
 a2111o_1 _20720_ (.A1(net1091),
    .A2(_05516_),
    .B1(_05518_),
    .C1(_05519_),
    .D1(_05521_),
    .X(_05522_));
 a21oi_1 _20721_ (.A1(_05514_),
    .A2(_05522_),
    .B1(net1097),
    .Y(_05523_));
 o32a_1 _20722_ (.A1(_07832_),
    .A2(_05511_),
    .A3(_05523_),
    .B1(_05512_),
    .B2(net1322),
    .X(_01261_));
 nor2_1 _20723_ (.A(_07827_),
    .B(_10718_),
    .Y(_05524_));
 or2_1 _20724_ (.A(\digitop_pav2.boot_inst.boot_ctrl0.proc_boot_end_i ),
    .B(_05524_),
    .X(_01262_));
 nand3_1 _20725_ (.A(\digitop_pav2.boot_inst.boot_proc0.proc_stage[0] ),
    .B(net1325),
    .C(_07833_),
    .Y(_05525_));
 mux2_1 _20726_ (.A0(net1134),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[16] ),
    .S(net1308),
    .X(_01263_));
 mux2_1 _20727_ (.A0(net1131),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[17] ),
    .S(net1308),
    .X(_01264_));
 mux2_1 _20728_ (.A0(net1127),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[18] ),
    .S(net1307),
    .X(_01265_));
 mux2_1 _20729_ (.A0(net1124),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[19] ),
    .S(net1307),
    .X(_01266_));
 mux2_1 _20730_ (.A0(net1121),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[20] ),
    .S(net1307),
    .X(_01267_));
 mux2_1 _20731_ (.A0(net1119),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[21] ),
    .S(net1307),
    .X(_01268_));
 mux2_1 _20732_ (.A0(net1116),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[22] ),
    .S(net1307),
    .X(_01269_));
 mux2_1 _20733_ (.A0(net1111),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[23] ),
    .S(net1307),
    .X(_01270_));
 mux2_1 _20734_ (.A0(net1109),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[24] ),
    .S(net1307),
    .X(_01271_));
 mux2_1 _20735_ (.A0(net1104),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[25] ),
    .S(net1308),
    .X(_01272_));
 mux2_1 _20736_ (.A0(net1101),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[26] ),
    .S(net1308),
    .X(_01273_));
 mux2_1 _20737_ (.A0(net1097),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[27] ),
    .S(net1308),
    .X(_01274_));
 mux2_1 _20738_ (.A0(net1095),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[28] ),
    .S(net1308),
    .X(_01275_));
 mux2_1 _20739_ (.A0(net1091),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[29] ),
    .S(net1307),
    .X(_01276_));
 mux2_1 _20740_ (.A0(net1088),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[30] ),
    .S(net1307),
    .X(_01277_));
 mux2_1 _20741_ (.A0(net1085),
    .A1(\digitop_pav2.boot_inst.boot_proc0.proc_mask[31] ),
    .S(net1307),
    .X(_01278_));
 a22o_1 _20742_ (.A1(\digitop_pav2.boot_inst.boot_ctrl0.replay ),
    .A2(net1400),
    .B1(_07829_),
    .B2(_07831_),
    .X(_01279_));
 mux2_1 _20743_ (.A0(\digitop_pav2.boot_inst.boot_proc0.proc_boot_sync ),
    .A1(\digitop_pav2.boot_inst.boot_ctrl0.proc_boot_end_i ),
    .S(_05524_),
    .X(_01280_));
 a31o_1 _20744_ (.A1(\digitop_pav2.boot_inst.boot_proc0.proc_boot_sync ),
    .A2(_07837_),
    .A3(_05524_),
    .B1(\digitop_pav2.boot_inst.boot_ctrl0.proc_crc_end_i ),
    .X(_01281_));
 nand2_1 _20745_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_0.A ),
    .B(_07518_),
    .Y(_05526_));
 or2_1 _20746_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_0.A ),
    .B(_07518_),
    .X(_05527_));
 nand2_1 _20747_ (.A(_05526_),
    .B(_05527_),
    .Y(_05528_));
 mux2_1 _20748_ (.A0(_05528_),
    .A1(_10797_),
    .S(_10799_),
    .X(_05529_));
 inv_2 _20749_ (.A(_05529_),
    .Y(_01282_));
 xnor2_1 _20750_ (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_0.A ),
    .B(_05526_),
    .Y(_05530_));
 mux2_1 _20751_ (.A0(_05530_),
    .A1(_10793_),
    .S(_10799_),
    .X(_01283_));
 nand2_4 _20752_ (.A(net468),
    .B(net173),
    .Y(_05531_));
 and4b_4 _20753_ (.A_N(_11194_),
    .B(_02735_),
    .C(_03427_),
    .D(_05531_),
    .X(_05532_));
 nand4b_4 _20754_ (.A_N(_11194_),
    .B(_02735_),
    .C(_03427_),
    .D(_05531_),
    .Y(_05533_));
 xor2_1 _20755_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[0] ),
    .X(_05534_));
 o21ai_1 _20756_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[0] ),
    .B1(net433),
    .Y(_05535_));
 a21oi_1 _20757_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[0] ),
    .B1(_05535_),
    .Y(_05536_));
 a211o_1 _20758_ (.A1(net419),
    .A2(_05534_),
    .B1(_05536_),
    .C1(_05533_),
    .X(_05537_));
 o32a_1 _20759_ (.A1(_11393_),
    .A2(_02747_),
    .A3(_05537_),
    .B1(_05532_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[0] ),
    .X(_01288_));
 o21ai_1 _20760_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[1] ),
    .B1(net432),
    .Y(_05538_));
 a21oi_1 _20761_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[1] ),
    .B1(_05538_),
    .Y(_05539_));
 xor2_1 _20762_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[1] ),
    .X(_05540_));
 a211o_1 _20763_ (.A1(net420),
    .A2(_05540_),
    .B1(_05539_),
    .C1(_05533_),
    .X(_05541_));
 o32a_1 _20764_ (.A1(_02182_),
    .A2(_02758_),
    .A3(_05541_),
    .B1(_05532_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[1] ),
    .X(_01289_));
 o21ai_1 _20765_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[2] ),
    .B1(net435),
    .Y(_05542_));
 a21oi_1 _20766_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[2] ),
    .B1(_05542_),
    .Y(_05543_));
 xor2_1 _20767_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[2] ),
    .X(_05544_));
 a2111o_1 _20768_ (.A1(net421),
    .A2(_05544_),
    .B1(_05543_),
    .C1(_05533_),
    .D1(_02280_),
    .X(_05545_));
 o32a_1 _20769_ (.A1(_02265_),
    .A2(_02767_),
    .A3(_05545_),
    .B1(_05532_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[2] ),
    .X(_01290_));
 or2_1 _20770_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[3] ),
    .X(_05546_));
 nand2_1 _20771_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[3] ),
    .Y(_05547_));
 or2_1 _20772_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[3] ),
    .X(_05548_));
 nand2_1 _20773_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state5_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[3] ),
    .Y(_05549_));
 a311o_1 _20774_ (.A1(net436),
    .A2(_05548_),
    .A3(_05549_),
    .B1(_02354_),
    .C1(_05533_),
    .X(_05550_));
 a31o_1 _20775_ (.A1(net422),
    .A2(_05546_),
    .A3(_05547_),
    .B1(_05550_),
    .X(_05551_));
 o32a_1 _20776_ (.A1(_02339_),
    .A2(_02779_),
    .A3(_05551_),
    .B1(_05532_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[3] ),
    .X(_01291_));
 xor2_1 _20777_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[4] ),
    .X(_05552_));
 o21ai_1 _20778_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[4] ),
    .B1(net436),
    .Y(_05553_));
 a21oi_1 _20779_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[4] ),
    .B1(_05553_),
    .Y(_05554_));
 a2111o_1 _20780_ (.A1(net422),
    .A2(_05552_),
    .B1(_05554_),
    .C1(_02423_),
    .D1(_05533_),
    .X(_05555_));
 o32a_1 _20781_ (.A1(_02413_),
    .A2(_02788_),
    .A3(_05555_),
    .B1(_05532_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[4] ),
    .X(_01292_));
 or2_1 _20782_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[5] ),
    .X(_05556_));
 nand2_1 _20783_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[5] ),
    .Y(_05557_));
 o21ai_1 _20784_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[5] ),
    .B1(net437),
    .Y(_05558_));
 a21oi_1 _20785_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[5] ),
    .B1(_05558_),
    .Y(_05559_));
 a31o_1 _20786_ (.A1(net423),
    .A2(_05556_),
    .A3(_05557_),
    .B1(_05559_),
    .X(_05560_));
 or4_1 _20787_ (.A(_02511_),
    .B(_02794_),
    .C(_05533_),
    .D(_05560_),
    .X(_05561_));
 o22a_1 _20788_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[5] ),
    .A2(_05532_),
    .B1(_05561_),
    .B2(_02482_),
    .X(_01293_));
 o21ai_1 _20789_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[6] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[6] ),
    .B1(net432),
    .Y(_05562_));
 a21oi_1 _20790_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[6] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[6] ),
    .B1(_05562_),
    .Y(_05563_));
 xor2_1 _20791_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[6] ),
    .X(_05564_));
 a2111o_1 _20792_ (.A1(net418),
    .A2(_05564_),
    .B1(_05563_),
    .C1(_05533_),
    .D1(_02562_),
    .X(_05565_));
 o32a_1 _20793_ (.A1(_02552_),
    .A2(_02811_),
    .A3(_05565_),
    .B1(_05532_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state5_r[6] ),
    .X(_01294_));
 or2_1 _20794_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[7] ),
    .X(_05566_));
 nand2_1 _20795_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[7] ),
    .Y(_05567_));
 o21ai_1 _20796_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[7] ),
    .B1(net430),
    .Y(_05568_));
 a21oi_1 _20797_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key5_r[7] ),
    .B1(_05568_),
    .Y(_05569_));
 a311o_1 _20798_ (.A1(net415),
    .A2(_05566_),
    .A3(_05567_),
    .B1(_05569_),
    .C1(_05533_),
    .X(_05570_));
 o22a_1 _20799_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ),
    .A2(_05532_),
    .B1(_05570_),
    .B2(_03614_),
    .X(_01295_));
 nor2_1 _20800_ (.A(_11216_),
    .B(net343),
    .Y(_05571_));
 or2_2 _20801_ (.A(_11216_),
    .B(net343),
    .X(_05572_));
 nand2_1 _20802_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[0] ),
    .Y(_05573_));
 or2_1 _20803_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[0] ),
    .X(_05574_));
 a31o_1 _20804_ (.A1(net454),
    .A2(_05573_),
    .A3(_05574_),
    .B1(net318),
    .X(_05575_));
 o22a_1 _20805_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[0] ),
    .A2(net320),
    .B1(_05575_),
    .B2(_05442_),
    .X(_01296_));
 nand2_1 _20806_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[1] ),
    .Y(_05576_));
 or2_1 _20807_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[1] ),
    .X(_05577_));
 a31o_1 _20808_ (.A1(net454),
    .A2(_05576_),
    .A3(_05577_),
    .B1(net319),
    .X(_05578_));
 o22a_1 _20809_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[1] ),
    .A2(net321),
    .B1(_05578_),
    .B2(_05446_),
    .X(_01297_));
 or2_1 _20810_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[2] ),
    .X(_05579_));
 nand2_1 _20811_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[2] ),
    .Y(_05580_));
 a31o_1 _20812_ (.A1(net451),
    .A2(_05579_),
    .A3(_05580_),
    .B1(net319),
    .X(_05581_));
 o22a_1 _20813_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[2] ),
    .A2(net321),
    .B1(_05581_),
    .B2(_05451_),
    .X(_01298_));
 nand2_1 _20814_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[3] ),
    .Y(_05582_));
 or2_1 _20815_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[3] ),
    .X(_05583_));
 a31o_1 _20816_ (.A1(net456),
    .A2(_05582_),
    .A3(_05583_),
    .B1(net319),
    .X(_05584_));
 o22a_1 _20817_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[3] ),
    .A2(net321),
    .B1(_05584_),
    .B2(_05456_),
    .X(_01299_));
 or2_1 _20818_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[4] ),
    .X(_05585_));
 nand2_1 _20819_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[4] ),
    .Y(_05586_));
 a31o_1 _20820_ (.A1(net457),
    .A2(_05585_),
    .A3(_05586_),
    .B1(net319),
    .X(_05587_));
 o22a_1 _20821_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[4] ),
    .A2(net321),
    .B1(_05587_),
    .B2(_05460_),
    .X(_01300_));
 or2_1 _20822_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[5] ),
    .X(_05588_));
 nand2_1 _20823_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[5] ),
    .Y(_05589_));
 a31o_1 _20824_ (.A1(net465),
    .A2(_05588_),
    .A3(_05589_),
    .B1(net319),
    .X(_05590_));
 o22a_1 _20825_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[5] ),
    .A2(net321),
    .B1(_05590_),
    .B2(_05465_),
    .X(_01301_));
 nand2_1 _20826_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[6] ),
    .Y(_05591_));
 or2_1 _20827_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[6] ),
    .X(_05592_));
 a31o_1 _20828_ (.A1(net454),
    .A2(_05591_),
    .A3(_05592_),
    .B1(net319),
    .X(_05593_));
 o22a_1 _20829_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[6] ),
    .A2(net321),
    .B1(_05593_),
    .B2(_05470_),
    .X(_01302_));
 or2_1 _20830_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[7] ),
    .X(_05594_));
 nand2_1 _20831_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[7] ),
    .Y(_05595_));
 a31o_1 _20832_ (.A1(net459),
    .A2(_05594_),
    .A3(_05595_),
    .B1(net318),
    .X(_05596_));
 o22a_1 _20833_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[7] ),
    .A2(net320),
    .B1(_05596_),
    .B2(_05473_),
    .X(_01303_));
 or2_1 _20834_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[8] ),
    .X(_05597_));
 nand2_1 _20835_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[8] ),
    .Y(_05598_));
 a31o_1 _20836_ (.A1(net461),
    .A2(_05597_),
    .A3(_05598_),
    .B1(net318),
    .X(_05599_));
 o22a_1 _20837_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[8] ),
    .A2(net320),
    .B1(_05599_),
    .B2(_05477_),
    .X(_01304_));
 nand2_1 _20838_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[9] ),
    .Y(_05600_));
 or2_1 _20839_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[9] ),
    .X(_05601_));
 a31o_1 _20840_ (.A1(net442),
    .A2(_05600_),
    .A3(_05601_),
    .B1(net318),
    .X(_05602_));
 o22a_1 _20841_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[9] ),
    .A2(net320),
    .B1(_05602_),
    .B2(_05480_),
    .X(_01305_));
 nand2_1 _20842_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[10] ),
    .Y(_05603_));
 or2_1 _20843_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[10] ),
    .X(_05604_));
 a31o_1 _20844_ (.A1(net447),
    .A2(_05603_),
    .A3(_05604_),
    .B1(net318),
    .X(_05605_));
 o22a_1 _20845_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[10] ),
    .A2(net320),
    .B1(_05605_),
    .B2(_05484_),
    .X(_01306_));
 nand2_1 _20846_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[11] ),
    .Y(_05606_));
 or2_1 _20847_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[11] ),
    .X(_05607_));
 a31o_1 _20848_ (.A1(net461),
    .A2(_05606_),
    .A3(_05607_),
    .B1(net318),
    .X(_05608_));
 o22a_1 _20849_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[11] ),
    .A2(net320),
    .B1(_05608_),
    .B2(_05489_),
    .X(_01307_));
 nand2_1 _20850_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[12] ),
    .Y(_05609_));
 or2_1 _20851_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[12] ),
    .X(_05610_));
 a31o_1 _20852_ (.A1(net461),
    .A2(_05609_),
    .A3(_05610_),
    .B1(net318),
    .X(_05611_));
 o22a_1 _20853_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[12] ),
    .A2(net320),
    .B1(_05611_),
    .B2(_05494_),
    .X(_01308_));
 nand2_1 _20854_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[13] ),
    .Y(_05612_));
 or2_1 _20855_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[13] ),
    .X(_05613_));
 a31o_1 _20856_ (.A1(net462),
    .A2(_05612_),
    .A3(_05613_),
    .B1(net318),
    .X(_05614_));
 o22a_1 _20857_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[13] ),
    .A2(net320),
    .B1(_05614_),
    .B2(_05499_),
    .X(_01309_));
 nand2_1 _20858_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[14] ),
    .Y(_05615_));
 or2_1 _20859_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[14] ),
    .X(_05616_));
 a31o_1 _20860_ (.A1(net443),
    .A2(_05615_),
    .A3(_05616_),
    .B1(net318),
    .X(_05617_));
 o22a_1 _20861_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[14] ),
    .A2(net320),
    .B1(_05617_),
    .B2(_05504_),
    .X(_01310_));
 nand2_1 _20862_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[15] ),
    .Y(_05618_));
 or2_1 _20863_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[15] ),
    .X(_05619_));
 a31o_1 _20864_ (.A1(net442),
    .A2(_05618_),
    .A3(_05619_),
    .B1(net318),
    .X(_05620_));
 o22a_1 _20865_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key4_r[15] ),
    .A2(net320),
    .B1(_05620_),
    .B2(_05507_),
    .X(_01311_));
 nor2_2 _20866_ (.A(_11202_),
    .B(net343),
    .Y(_05621_));
 or2_2 _20867_ (.A(_11202_),
    .B(net344),
    .X(_05622_));
 or2_1 _20868_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[0] ),
    .X(_05623_));
 nand2_1 _20869_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[0] ),
    .Y(_05624_));
 a31o_1 _20870_ (.A1(net454),
    .A2(_05623_),
    .A3(_05624_),
    .B1(net314),
    .X(_05625_));
 o22a_1 _20871_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[0] ),
    .A2(net316),
    .B1(_05625_),
    .B2(_05442_),
    .X(_01312_));
 nand2_1 _20872_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[1] ),
    .Y(_05626_));
 or2_1 _20873_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[1] ),
    .X(_05627_));
 a31o_1 _20874_ (.A1(net453),
    .A2(_05626_),
    .A3(_05627_),
    .B1(net315),
    .X(_05628_));
 o22a_1 _20875_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[1] ),
    .A2(net317),
    .B1(_05628_),
    .B2(_05446_),
    .X(_01313_));
 nand2_1 _20876_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[2] ),
    .Y(_05629_));
 or2_1 _20877_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[2] ),
    .X(_05630_));
 a31o_1 _20878_ (.A1(net451),
    .A2(_05629_),
    .A3(_05630_),
    .B1(net315),
    .X(_05631_));
 o22a_1 _20879_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[2] ),
    .A2(net317),
    .B1(_05631_),
    .B2(_05451_),
    .X(_01314_));
 nand2_1 _20880_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[3] ),
    .Y(_05632_));
 or2_1 _20881_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[3] ),
    .X(_05633_));
 a31o_1 _20882_ (.A1(net455),
    .A2(_05632_),
    .A3(_05633_),
    .B1(net315),
    .X(_05634_));
 o22a_1 _20883_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[3] ),
    .A2(net317),
    .B1(_05634_),
    .B2(_05456_),
    .X(_01315_));
 or2_1 _20884_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[4] ),
    .X(_05635_));
 nand2_1 _20885_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[4] ),
    .Y(_05636_));
 a31o_1 _20886_ (.A1(net457),
    .A2(_05635_),
    .A3(_05636_),
    .B1(net315),
    .X(_05637_));
 o22a_1 _20887_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[4] ),
    .A2(net317),
    .B1(_05637_),
    .B2(_05460_),
    .X(_01316_));
 or2_1 _20888_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[5] ),
    .X(_05638_));
 nand2_1 _20889_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[5] ),
    .Y(_05639_));
 a31o_1 _20890_ (.A1(net457),
    .A2(_05638_),
    .A3(_05639_),
    .B1(net315),
    .X(_05640_));
 o22a_1 _20891_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[5] ),
    .A2(net317),
    .B1(_05640_),
    .B2(_05465_),
    .X(_01317_));
 nand2_1 _20892_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[6] ),
    .Y(_05641_));
 or2_1 _20893_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[6] ),
    .X(_05642_));
 a31o_1 _20894_ (.A1(net452),
    .A2(_05641_),
    .A3(_05642_),
    .B1(net315),
    .X(_05643_));
 o22a_1 _20895_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[6] ),
    .A2(net317),
    .B1(_05643_),
    .B2(_05470_),
    .X(_01318_));
 or2_1 _20896_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[7] ),
    .X(_05644_));
 nand2_1 _20897_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key5_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[7] ),
    .Y(_05645_));
 a31o_1 _20898_ (.A1(net444),
    .A2(_05644_),
    .A3(_05645_),
    .B1(net314),
    .X(_05646_));
 o22a_1 _20899_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[7] ),
    .A2(net316),
    .B1(_05646_),
    .B2(_05473_),
    .X(_01319_));
 or2_1 _20900_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[8] ),
    .X(_05647_));
 nand2_1 _20901_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[8] ),
    .Y(_05648_));
 a31o_1 _20902_ (.A1(net460),
    .A2(_05647_),
    .A3(_05648_),
    .B1(net314),
    .X(_05649_));
 o22a_1 _20903_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[8] ),
    .A2(net316),
    .B1(_05649_),
    .B2(_05477_),
    .X(_01320_));
 nand2_1 _20904_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[9] ),
    .Y(_05650_));
 or2_1 _20905_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[9] ),
    .X(_05651_));
 a31o_1 _20906_ (.A1(net443),
    .A2(_05650_),
    .A3(_05651_),
    .B1(net314),
    .X(_05652_));
 o22a_1 _20907_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[9] ),
    .A2(net316),
    .B1(_05652_),
    .B2(_05480_),
    .X(_01321_));
 nand2_1 _20908_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[10] ),
    .Y(_05653_));
 or2_1 _20909_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[10] ),
    .X(_05654_));
 a31o_1 _20910_ (.A1(net448),
    .A2(_05653_),
    .A3(_05654_),
    .B1(net314),
    .X(_05655_));
 o22a_1 _20911_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[10] ),
    .A2(net316),
    .B1(_05655_),
    .B2(_05484_),
    .X(_01322_));
 nand2_1 _20912_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[11] ),
    .Y(_05656_));
 or2_1 _20913_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[11] ),
    .X(_05657_));
 a31o_1 _20914_ (.A1(net460),
    .A2(_05656_),
    .A3(_05657_),
    .B1(net314),
    .X(_05658_));
 o22a_1 _20915_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[11] ),
    .A2(net316),
    .B1(_05658_),
    .B2(_05489_),
    .X(_01323_));
 nand2_1 _20916_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[12] ),
    .Y(_05659_));
 or2_1 _20917_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[12] ),
    .X(_05660_));
 a31o_1 _20918_ (.A1(net461),
    .A2(_05659_),
    .A3(_05660_),
    .B1(net314),
    .X(_05661_));
 o22a_1 _20919_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[12] ),
    .A2(net316),
    .B1(_05661_),
    .B2(_05494_),
    .X(_01324_));
 nand2_1 _20920_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[13] ),
    .Y(_05662_));
 or2_1 _20921_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[13] ),
    .X(_05663_));
 a31o_1 _20922_ (.A1(net462),
    .A2(_05662_),
    .A3(_05663_),
    .B1(net314),
    .X(_05664_));
 o22a_1 _20923_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[13] ),
    .A2(net316),
    .B1(_05664_),
    .B2(_05499_),
    .X(_01325_));
 nand2_1 _20924_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[14] ),
    .Y(_05665_));
 or2_1 _20925_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[14] ),
    .X(_05666_));
 a31o_1 _20926_ (.A1(net448),
    .A2(_05665_),
    .A3(_05666_),
    .B1(net314),
    .X(_05667_));
 o22a_1 _20927_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[14] ),
    .A2(net316),
    .B1(_05667_),
    .B2(_05504_),
    .X(_01326_));
 nand2_1 _20928_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[15] ),
    .Y(_05668_));
 or2_1 _20929_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key3_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key5_r[15] ),
    .X(_05669_));
 a31o_1 _20930_ (.A1(net448),
    .A2(_05668_),
    .A3(_05669_),
    .B1(net314),
    .X(_05670_));
 o22a_1 _20931_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key3_r[15] ),
    .A2(net316),
    .B1(_05670_),
    .B2(_05507_),
    .X(_01327_));
 and2_1 _20932_ (.A(net365),
    .B(_05435_),
    .X(_05671_));
 o21ai_1 _20933_ (.A1(net409),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[0] ),
    .B1(net299),
    .Y(_05672_));
 a31o_1 _20934_ (.A1(net455),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[0] ),
    .A3(_07227_),
    .B1(_05442_),
    .X(_05673_));
 a22o_1 _20935_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[0] ),
    .A2(_05672_),
    .B1(_05673_),
    .B2(net299),
    .X(_01328_));
 o21ai_1 _20936_ (.A1(net408),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[1] ),
    .B1(net299),
    .Y(_05674_));
 a31o_1 _20937_ (.A1(net454),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[1] ),
    .A3(_07228_),
    .B1(_05446_),
    .X(_05675_));
 a22o_1 _20938_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[1] ),
    .A2(_05674_),
    .B1(_05675_),
    .B2(net299),
    .X(_01329_));
 o21ai_1 _20939_ (.A1(net407),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[2] ),
    .B1(net299),
    .Y(_05676_));
 a31o_1 _20940_ (.A1(net450),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[2] ),
    .A3(_07229_),
    .B1(_05451_),
    .X(_05677_));
 a22o_1 _20941_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[2] ),
    .A2(_05676_),
    .B1(_05677_),
    .B2(net299),
    .X(_01330_));
 o21ai_1 _20942_ (.A1(net409),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[3] ),
    .B1(net300),
    .Y(_05678_));
 a31o_1 _20943_ (.A1(net455),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[3] ),
    .A3(_07230_),
    .B1(_05456_),
    .X(_05679_));
 a22o_1 _20944_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[3] ),
    .A2(_05678_),
    .B1(_05679_),
    .B2(net300),
    .X(_01331_));
 o21ai_1 _20945_ (.A1(net412),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[4] ),
    .B1(net299),
    .Y(_05680_));
 a31o_1 _20946_ (.A1(net465),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[4] ),
    .A3(_07231_),
    .B1(_05460_),
    .X(_05681_));
 a22o_1 _20947_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[4] ),
    .A2(_05680_),
    .B1(_05681_),
    .B2(net299),
    .X(_01332_));
 o21ai_1 _20948_ (.A1(net412),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[5] ),
    .B1(net300),
    .Y(_05682_));
 a31o_1 _20949_ (.A1(net465),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[5] ),
    .A3(_07232_),
    .B1(_05465_),
    .X(_05683_));
 a22o_1 _20950_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[5] ),
    .A2(_05682_),
    .B1(_05683_),
    .B2(net300),
    .X(_01333_));
 o21ai_1 _20951_ (.A1(net408),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[6] ),
    .B1(net299),
    .Y(_05684_));
 a31o_1 _20952_ (.A1(net451),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[6] ),
    .A3(_07233_),
    .B1(_05470_),
    .X(_05685_));
 a22o_1 _20953_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[6] ),
    .A2(_05684_),
    .B1(_05685_),
    .B2(net299),
    .X(_01334_));
 o21ai_1 _20954_ (.A1(net405),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[7] ),
    .B1(net297),
    .Y(_05686_));
 a31o_1 _20955_ (.A1(net445),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[7] ),
    .A3(_07234_),
    .B1(_05473_),
    .X(_05687_));
 a22o_1 _20956_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[7] ),
    .A2(_05686_),
    .B1(_05687_),
    .B2(net297),
    .X(_01335_));
 o21ai_1 _20957_ (.A1(net410),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[8] ),
    .B1(net298),
    .Y(_05688_));
 a31o_1 _20958_ (.A1(net448),
    .A2(_07171_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key4_r[8] ),
    .B1(_05477_),
    .X(_05689_));
 a22o_1 _20959_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[8] ),
    .A2(_05688_),
    .B1(_05689_),
    .B2(net298),
    .X(_01336_));
 o21ai_1 _20960_ (.A1(net405),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[9] ),
    .B1(net297),
    .Y(_05690_));
 a31o_1 _20961_ (.A1(net443),
    .A2(_07173_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key4_r[9] ),
    .B1(_05480_),
    .X(_05691_));
 a22o_1 _20962_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[9] ),
    .A2(_05690_),
    .B1(_05691_),
    .B2(net297),
    .X(_01337_));
 o21ai_1 _20963_ (.A1(net406),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[10] ),
    .B1(net297),
    .Y(_05692_));
 a31o_1 _20964_ (.A1(net447),
    .A2(_07175_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key4_r[10] ),
    .B1(_05484_),
    .X(_05693_));
 a22o_1 _20965_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[10] ),
    .A2(_05692_),
    .B1(_05693_),
    .B2(net297),
    .X(_01338_));
 o21ai_1 _20966_ (.A1(net410),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[11] ),
    .B1(net298),
    .Y(_05694_));
 a31o_1 _20967_ (.A1(net460),
    .A2(_07177_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key4_r[11] ),
    .B1(_05489_),
    .X(_05695_));
 a22o_1 _20968_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[11] ),
    .A2(_05694_),
    .B1(_05695_),
    .B2(net298),
    .X(_01339_));
 o21ai_1 _20969_ (.A1(net410),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[12] ),
    .B1(net298),
    .Y(_05696_));
 a31o_1 _20970_ (.A1(net460),
    .A2(_07179_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key4_r[12] ),
    .B1(_05494_),
    .X(_05697_));
 a22o_1 _20971_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[12] ),
    .A2(_05696_),
    .B1(_05697_),
    .B2(net298),
    .X(_01340_));
 o21ai_1 _20972_ (.A1(net410),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[13] ),
    .B1(net298),
    .Y(_05698_));
 a31o_1 _20973_ (.A1(net462),
    .A2(_07181_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key4_r[13] ),
    .B1(_05499_),
    .X(_05699_));
 a22o_1 _20974_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[13] ),
    .A2(_05698_),
    .B1(_05699_),
    .B2(net298),
    .X(_01341_));
 o21ai_1 _20975_ (.A1(net405),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[14] ),
    .B1(net297),
    .Y(_05700_));
 a31o_1 _20976_ (.A1(net443),
    .A2(_07183_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key4_r[14] ),
    .B1(_05504_),
    .X(_05701_));
 a22o_1 _20977_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[14] ),
    .A2(_05700_),
    .B1(_05701_),
    .B2(net297),
    .X(_01342_));
 o21ai_1 _20978_ (.A1(net406),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[15] ),
    .B1(net297),
    .Y(_05702_));
 a31o_1 _20979_ (.A1(net442),
    .A2(_07185_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key4_r[15] ),
    .B1(_05507_),
    .X(_05703_));
 a22o_1 _20980_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key2_r[15] ),
    .A2(_05702_),
    .B1(_05703_),
    .B2(net297),
    .X(_01343_));
 and2_1 _20981_ (.A(net355),
    .B(_05435_),
    .X(_05704_));
 o21ai_1 _20982_ (.A1(net408),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[0] ),
    .B1(net295),
    .Y(_05705_));
 a31o_1 _20983_ (.A1(net454),
    .A2(_07198_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[0] ),
    .B1(_05442_),
    .X(_05706_));
 a22o_1 _20984_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[0] ),
    .A2(_05705_),
    .B1(_05706_),
    .B2(net295),
    .X(_01344_));
 o21ai_1 _20985_ (.A1(net408),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[1] ),
    .B1(net295),
    .Y(_05707_));
 a31o_1 _20986_ (.A1(net453),
    .A2(_07196_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[1] ),
    .B1(_05446_),
    .X(_05708_));
 a22o_1 _20987_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[1] ),
    .A2(_05707_),
    .B1(_05708_),
    .B2(net295),
    .X(_01345_));
 o21ai_1 _20988_ (.A1(net407),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[2] ),
    .B1(net295),
    .Y(_05709_));
 a31o_1 _20989_ (.A1(net450),
    .A2(_07200_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[2] ),
    .B1(_05451_),
    .X(_05710_));
 a22o_1 _20990_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[2] ),
    .A2(_05709_),
    .B1(_05710_),
    .B2(net295),
    .X(_01346_));
 o21ai_1 _20991_ (.A1(net409),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[3] ),
    .B1(net295),
    .Y(_05711_));
 a31o_1 _20992_ (.A1(net455),
    .A2(_07202_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[3] ),
    .B1(_05456_),
    .X(_05712_));
 a22o_1 _20993_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[3] ),
    .A2(_05711_),
    .B1(_05712_),
    .B2(net295),
    .X(_01347_));
 o21ai_1 _20994_ (.A1(net409),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[4] ),
    .B1(net296),
    .Y(_05713_));
 a31o_1 _20995_ (.A1(net457),
    .A2(_07204_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[4] ),
    .B1(_05460_),
    .X(_05714_));
 a22o_1 _20996_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[4] ),
    .A2(_05713_),
    .B1(_05714_),
    .B2(net296),
    .X(_01348_));
 o21ai_1 _20997_ (.A1(net412),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[5] ),
    .B1(net296),
    .Y(_05715_));
 a31o_1 _20998_ (.A1(net457),
    .A2(_07206_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[5] ),
    .B1(_05465_),
    .X(_05716_));
 a22o_1 _20999_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[5] ),
    .A2(_05715_),
    .B1(_05716_),
    .B2(net296),
    .X(_01349_));
 o21ai_1 _21000_ (.A1(net407),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[6] ),
    .B1(net295),
    .Y(_05717_));
 a31o_1 _21001_ (.A1(net451),
    .A2(_07208_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[6] ),
    .B1(_05470_),
    .X(_05718_));
 a22o_1 _21002_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[6] ),
    .A2(_05717_),
    .B1(_05718_),
    .B2(net295),
    .X(_01350_));
 o21ai_1 _21003_ (.A1(net405),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[7] ),
    .B1(net294),
    .Y(_05719_));
 a31o_1 _21004_ (.A1(net444),
    .A2(_07210_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[7] ),
    .B1(_05473_),
    .X(_05720_));
 a22o_1 _21005_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[7] ),
    .A2(_05719_),
    .B1(_05720_),
    .B2(net294),
    .X(_01351_));
 o21ai_1 _21006_ (.A1(net410),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[8] ),
    .B1(net292),
    .Y(_05721_));
 a31o_1 _21007_ (.A1(net447),
    .A2(_07187_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[8] ),
    .B1(_05477_),
    .X(_05722_));
 a22o_1 _21008_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[8] ),
    .A2(_05721_),
    .B1(_05722_),
    .B2(net292),
    .X(_01352_));
 o21ai_1 _21009_ (.A1(net405),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[9] ),
    .B1(net294),
    .Y(_05723_));
 a31o_1 _21010_ (.A1(net446),
    .A2(_07188_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[9] ),
    .B1(_05480_),
    .X(_05724_));
 a22o_1 _21011_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[9] ),
    .A2(_05723_),
    .B1(_05724_),
    .B2(net294),
    .X(_01353_));
 o21ai_1 _21012_ (.A1(net406),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[10] ),
    .B1(net292),
    .Y(_05725_));
 a31o_1 _21013_ (.A1(net447),
    .A2(_07189_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[10] ),
    .B1(_05484_),
    .X(_05726_));
 a22o_1 _21014_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[10] ),
    .A2(_05725_),
    .B1(_05726_),
    .B2(net292),
    .X(_01354_));
 o21ai_1 _21015_ (.A1(net410),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[11] ),
    .B1(net292),
    .Y(_05727_));
 a31o_1 _21016_ (.A1(net460),
    .A2(_07190_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[11] ),
    .B1(_05489_),
    .X(_05728_));
 a22o_1 _21017_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[11] ),
    .A2(_05727_),
    .B1(_05728_),
    .B2(net292),
    .X(_01355_));
 o21ai_1 _21018_ (.A1(net410),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[12] ),
    .B1(net293),
    .Y(_05729_));
 a31o_1 _21019_ (.A1(net460),
    .A2(_07191_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[12] ),
    .B1(_05494_),
    .X(_05730_));
 a22o_1 _21020_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[12] ),
    .A2(_05729_),
    .B1(_05730_),
    .B2(net293),
    .X(_01356_));
 o21ai_1 _21021_ (.A1(net410),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[13] ),
    .B1(net293),
    .Y(_05731_));
 a31o_1 _21022_ (.A1(net462),
    .A2(_07192_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[13] ),
    .B1(_05499_),
    .X(_05732_));
 a22o_1 _21023_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[13] ),
    .A2(_05731_),
    .B1(_05732_),
    .B2(net293),
    .X(_01357_));
 o21ai_1 _21024_ (.A1(net405),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[14] ),
    .B1(net292),
    .Y(_05733_));
 a31o_1 _21025_ (.A1(net448),
    .A2(_07193_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[14] ),
    .B1(_05504_),
    .X(_05734_));
 a22o_1 _21026_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[14] ),
    .A2(_05733_),
    .B1(_05734_),
    .B2(net292),
    .X(_01358_));
 o21ai_1 _21027_ (.A1(net406),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key3_r[15] ),
    .B1(net292),
    .Y(_05735_));
 a31o_1 _21028_ (.A1(net448),
    .A2(_07194_),
    .A3(\digitop_pav2.aes128_inst.aes128_regs.key3_r[15] ),
    .B1(_05507_),
    .X(_05736_));
 a22o_1 _21029_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key1_r[15] ),
    .A2(_05735_),
    .B1(_05736_),
    .B2(net292),
    .X(_01359_));
 nor2_1 _21030_ (.A(net393),
    .B(net345),
    .Y(_05737_));
 xor2_1 _21031_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[0] ),
    .B(_11392_),
    .X(_05738_));
 o21ai_1 _21032_ (.A1(net408),
    .A2(_05738_),
    .B1(net312),
    .Y(_05739_));
 o22a_1 _21033_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[0] ),
    .A2(net312),
    .B1(_05739_),
    .B2(_05442_),
    .X(_01360_));
 nand2_1 _21034_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[1] ),
    .B(_02181_),
    .Y(_05740_));
 or2_1 _21035_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[1] ),
    .B(_02181_),
    .X(_05741_));
 a311o_1 _21036_ (.A1(net453),
    .A2(_05740_),
    .A3(_05741_),
    .B1(net393),
    .C1(net345),
    .X(_05742_));
 o22a_1 _21037_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[1] ),
    .A2(net311),
    .B1(_05742_),
    .B2(_05446_),
    .X(_01361_));
 xor2_1 _21038_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[2] ),
    .B(_02264_),
    .X(_05743_));
 o21ai_1 _21039_ (.A1(net407),
    .A2(_05743_),
    .B1(net312),
    .Y(_05744_));
 o22a_1 _21040_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[2] ),
    .A2(net312),
    .B1(_05744_),
    .B2(_05451_),
    .X(_01362_));
 nand2_1 _21041_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[3] ),
    .B(_02338_),
    .Y(_05745_));
 or2_1 _21042_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[3] ),
    .B(_02338_),
    .X(_05746_));
 a311o_1 _21043_ (.A1(net455),
    .A2(_05745_),
    .A3(_05746_),
    .B1(net392),
    .C1(net345),
    .X(_05747_));
 o22a_1 _21044_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[3] ),
    .A2(net312),
    .B1(_05747_),
    .B2(_05456_),
    .X(_01363_));
 nand2_1 _21045_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[4] ),
    .B(_02412_),
    .Y(_05748_));
 or2_1 _21046_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[4] ),
    .B(_02412_),
    .X(_05749_));
 a311o_1 _21047_ (.A1(net458),
    .A2(_05748_),
    .A3(_05749_),
    .B1(net392),
    .C1(net345),
    .X(_05750_));
 o22a_1 _21048_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[4] ),
    .A2(net312),
    .B1(_05750_),
    .B2(_05460_),
    .X(_01364_));
 nand2_1 _21049_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[5] ),
    .B(net160),
    .Y(_05751_));
 or2_1 _21050_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[5] ),
    .B(net160),
    .X(_05752_));
 a311o_1 _21051_ (.A1(net457),
    .A2(_05751_),
    .A3(_05752_),
    .B1(net392),
    .C1(net346),
    .X(_05753_));
 o22a_1 _21052_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[5] ),
    .A2(net312),
    .B1(_05753_),
    .B2(_05465_),
    .X(_01365_));
 nand2_1 _21053_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[6] ),
    .B(_02551_),
    .Y(_05754_));
 or2_1 _21054_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[6] ),
    .B(_02551_),
    .X(_05755_));
 a311o_1 _21055_ (.A1(net452),
    .A2(_05754_),
    .A3(_05755_),
    .B1(net393),
    .C1(net345),
    .X(_05756_));
 o22a_1 _21056_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[6] ),
    .A2(net312),
    .B1(_05756_),
    .B2(_05470_),
    .X(_01366_));
 nand2_1 _21057_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[7] ),
    .B(_02615_),
    .Y(_05757_));
 or2_1 _21058_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[7] ),
    .B(_02615_),
    .X(_05758_));
 a311o_1 _21059_ (.A1(net446),
    .A2(_05757_),
    .A3(_05758_),
    .B1(net393),
    .C1(net343),
    .X(_05759_));
 o22a_1 _21060_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[7] ),
    .A2(net311),
    .B1(_05759_),
    .B2(_05473_),
    .X(_01367_));
 xor2_1 _21061_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[0] ),
    .X(_05760_));
 xnor2_1 _21062_ (.A(_02995_),
    .B(_05760_),
    .Y(_05761_));
 o21ai_1 _21063_ (.A1(net411),
    .A2(_05761_),
    .B1(net313),
    .Y(_05762_));
 o22a_1 _21064_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[8] ),
    .A2(net313),
    .B1(_05762_),
    .B2(_05477_),
    .X(_01368_));
 or2_1 _21065_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[1] ),
    .X(_05763_));
 nand2_1 _21066_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[1] ),
    .Y(_05764_));
 a21oi_1 _21067_ (.A1(_05763_),
    .A2(_05764_),
    .B1(_03081_),
    .Y(_05765_));
 a31o_1 _21068_ (.A1(_03081_),
    .A2(_05763_),
    .A3(_05764_),
    .B1(net405),
    .X(_05766_));
 o21ai_1 _21069_ (.A1(_05765_),
    .A2(_05766_),
    .B1(net311),
    .Y(_05767_));
 o22a_1 _21070_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[9] ),
    .A2(net311),
    .B1(_05767_),
    .B2(_05480_),
    .X(_01369_));
 xor2_1 _21071_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[2] ),
    .X(_05768_));
 xnor2_1 _21072_ (.A(_03149_),
    .B(_05768_),
    .Y(_05769_));
 o21ai_1 _21073_ (.A1(net406),
    .A2(_05769_),
    .B1(net311),
    .Y(_05770_));
 o22a_1 _21074_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[10] ),
    .A2(net311),
    .B1(_05770_),
    .B2(_05484_),
    .X(_01370_));
 or2_1 _21075_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[3] ),
    .X(_05771_));
 nand2_1 _21076_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[3] ),
    .Y(_05772_));
 a21oi_1 _21077_ (.A1(_05771_),
    .A2(_05772_),
    .B1(_03201_),
    .Y(_05773_));
 a31o_1 _21078_ (.A1(_03201_),
    .A2(_05771_),
    .A3(_05772_),
    .B1(net411),
    .X(_05774_));
 o21ai_1 _21079_ (.A1(_05773_),
    .A2(_05774_),
    .B1(net313),
    .Y(_05775_));
 o22a_1 _21080_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[11] ),
    .A2(net313),
    .B1(_05775_),
    .B2(_05489_),
    .X(_01371_));
 xor2_1 _21081_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[4] ),
    .X(_05776_));
 xnor2_1 _21082_ (.A(_03254_),
    .B(_05776_),
    .Y(_05777_));
 o21ai_1 _21083_ (.A1(net411),
    .A2(_05777_),
    .B1(net313),
    .Y(_05778_));
 o22a_1 _21084_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[12] ),
    .A2(net313),
    .B1(_05778_),
    .B2(_05494_),
    .X(_01372_));
 xor2_1 _21085_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[5] ),
    .X(_05779_));
 xnor2_1 _21086_ (.A(_03302_),
    .B(_05779_),
    .Y(_05780_));
 o21ai_1 _21087_ (.A1(net410),
    .A2(_05780_),
    .B1(net313),
    .Y(_05781_));
 o22a_1 _21088_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[13] ),
    .A2(net313),
    .B1(_05781_),
    .B2(_05499_),
    .X(_01373_));
 xor2_1 _21089_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[6] ),
    .X(_05782_));
 xnor2_1 _21090_ (.A(_03352_),
    .B(_05782_),
    .Y(_05783_));
 o21ai_1 _21091_ (.A1(net405),
    .A2(_05783_),
    .B1(net311),
    .Y(_05784_));
 o22a_1 _21092_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[14] ),
    .A2(net311),
    .B1(_05784_),
    .B2(_05504_),
    .X(_01374_));
 xor2_1 _21093_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key7_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[7] ),
    .X(_05785_));
 xnor2_1 _21094_ (.A(_03402_),
    .B(_05785_),
    .Y(_05786_));
 o21ai_1 _21095_ (.A1(net406),
    .A2(_05786_),
    .B1(net311),
    .Y(_05787_));
 o22a_1 _21096_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key7_r[15] ),
    .A2(net311),
    .B1(_05787_),
    .B2(_05507_),
    .X(_01375_));
 nor2_1 _21097_ (.A(net358),
    .B(net343),
    .Y(_05788_));
 xor2_1 _21098_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[0] ),
    .B(_11392_),
    .X(_05789_));
 o21ai_1 _21099_ (.A1(net408),
    .A2(_05789_),
    .B1(net310),
    .Y(_05790_));
 o22a_1 _21100_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[0] ),
    .A2(net310),
    .B1(_05790_),
    .B2(_05442_),
    .X(_01376_));
 nand2_1 _21101_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[1] ),
    .B(_02181_),
    .Y(_05791_));
 or2_1 _21102_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[1] ),
    .B(_02181_),
    .X(_05792_));
 a311o_1 _21103_ (.A1(net453),
    .A2(_05791_),
    .A3(_05792_),
    .B1(net359),
    .C1(net345),
    .X(_05793_));
 o22a_1 _21104_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[1] ),
    .A2(net310),
    .B1(_05793_),
    .B2(_05446_),
    .X(_01377_));
 xor2_1 _21105_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[2] ),
    .B(_02264_),
    .X(_05794_));
 o21ai_1 _21106_ (.A1(net407),
    .A2(_05794_),
    .B1(net310),
    .Y(_05795_));
 o22a_1 _21107_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[2] ),
    .A2(net310),
    .B1(_05795_),
    .B2(_05451_),
    .X(_01378_));
 nand2_1 _21108_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[3] ),
    .B(_02338_),
    .Y(_05796_));
 or2_1 _21109_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[3] ),
    .B(_02338_),
    .X(_05797_));
 a311o_1 _21110_ (.A1(net455),
    .A2(_05796_),
    .A3(_05797_),
    .B1(net359),
    .C1(net345),
    .X(_05798_));
 o22a_1 _21111_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[3] ),
    .A2(net310),
    .B1(_05798_),
    .B2(_05456_),
    .X(_01379_));
 nand2_1 _21112_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[4] ),
    .B(_02412_),
    .Y(_05799_));
 or2_1 _21113_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[4] ),
    .B(_02412_),
    .X(_05800_));
 a311o_1 _21114_ (.A1(net457),
    .A2(_05799_),
    .A3(_05800_),
    .B1(net359),
    .C1(net345),
    .X(_05801_));
 o22a_1 _21115_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[4] ),
    .A2(net309),
    .B1(_05801_),
    .B2(_05460_),
    .X(_01380_));
 nand2_1 _21116_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[5] ),
    .B(net160),
    .Y(_05802_));
 or2_1 _21117_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[5] ),
    .B(net160),
    .X(_05803_));
 a311o_1 _21118_ (.A1(net457),
    .A2(_05802_),
    .A3(_05803_),
    .B1(net359),
    .C1(net345),
    .X(_05804_));
 o22a_1 _21119_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[5] ),
    .A2(net310),
    .B1(_05804_),
    .B2(_05465_),
    .X(_01381_));
 nand2_1 _21120_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[6] ),
    .B(_02551_),
    .Y(_05805_));
 or2_1 _21121_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[6] ),
    .B(_02551_),
    .X(_05806_));
 a311o_1 _21122_ (.A1(net452),
    .A2(_05805_),
    .A3(_05806_),
    .B1(net359),
    .C1(net345),
    .X(_05807_));
 o22a_1 _21123_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[6] ),
    .A2(net310),
    .B1(_05807_),
    .B2(_05470_),
    .X(_01382_));
 nand2_1 _21124_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[7] ),
    .B(_02615_),
    .Y(_05808_));
 or2_1 _21125_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[7] ),
    .B(_02615_),
    .X(_05809_));
 a311o_1 _21126_ (.A1(net446),
    .A2(_05808_),
    .A3(_05809_),
    .B1(net358),
    .C1(net343),
    .X(_05810_));
 o22a_1 _21127_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[7] ),
    .A2(net309),
    .B1(_05810_),
    .B2(_05473_),
    .X(_01383_));
 nand2_1 _21128_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[8] ),
    .B(_02995_),
    .Y(_05811_));
 or2_1 _21129_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[8] ),
    .B(_02995_),
    .X(_05812_));
 a311o_1 _21130_ (.A1(net461),
    .A2(_05811_),
    .A3(_05812_),
    .B1(net358),
    .C1(net344),
    .X(_05813_));
 o22a_1 _21131_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[8] ),
    .A2(net309),
    .B1(_05813_),
    .B2(_05477_),
    .X(_01384_));
 nand2_1 _21132_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[9] ),
    .B(_03081_),
    .Y(_05814_));
 or2_1 _21133_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[9] ),
    .B(_03081_),
    .X(_05815_));
 a311o_1 _21134_ (.A1(net442),
    .A2(_05814_),
    .A3(_05815_),
    .B1(net358),
    .C1(net343),
    .X(_05816_));
 o22a_1 _21135_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[9] ),
    .A2(net309),
    .B1(_05816_),
    .B2(_05480_),
    .X(_01385_));
 nand2_1 _21136_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[10] ),
    .B(_03149_),
    .Y(_05817_));
 or2_1 _21137_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[10] ),
    .B(_03149_),
    .X(_05818_));
 a311o_1 _21138_ (.A1(net447),
    .A2(_05817_),
    .A3(_05818_),
    .B1(net358),
    .C1(net343),
    .X(_05819_));
 o22a_1 _21139_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[10] ),
    .A2(net309),
    .B1(_05819_),
    .B2(_05484_),
    .X(_01386_));
 or2_1 _21140_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[11] ),
    .B(_03201_),
    .X(_05820_));
 nand2_1 _21141_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[11] ),
    .B(_03201_),
    .Y(_05821_));
 a311o_1 _21142_ (.A1(net461),
    .A2(_05820_),
    .A3(_05821_),
    .B1(net359),
    .C1(net344),
    .X(_05822_));
 o22a_1 _21143_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[11] ),
    .A2(net309),
    .B1(_05822_),
    .B2(_05489_),
    .X(_01387_));
 nand2_1 _21144_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[12] ),
    .B(_03254_),
    .Y(_05823_));
 or2_1 _21145_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[12] ),
    .B(_03254_),
    .X(_05824_));
 a311o_1 _21146_ (.A1(net461),
    .A2(_05823_),
    .A3(_05824_),
    .B1(net358),
    .C1(net344),
    .X(_05825_));
 o22a_1 _21147_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[12] ),
    .A2(net309),
    .B1(_05825_),
    .B2(_05494_),
    .X(_01388_));
 nand2_1 _21148_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[13] ),
    .B(_03302_),
    .Y(_05826_));
 or2_1 _21149_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[13] ),
    .B(_03302_),
    .X(_05827_));
 a311o_1 _21150_ (.A1(net462),
    .A2(_05826_),
    .A3(_05827_),
    .B1(net358),
    .C1(net344),
    .X(_05828_));
 o22a_1 _21151_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[13] ),
    .A2(net309),
    .B1(_05828_),
    .B2(_05499_),
    .X(_01389_));
 nand2_1 _21152_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[14] ),
    .B(_03352_),
    .Y(_05829_));
 or2_1 _21153_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[14] ),
    .B(_03352_),
    .X(_05830_));
 a311o_1 _21154_ (.A1(net443),
    .A2(_05829_),
    .A3(_05830_),
    .B1(net358),
    .C1(net343),
    .X(_05831_));
 o22a_1 _21155_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[14] ),
    .A2(net309),
    .B1(_05831_),
    .B2(_05504_),
    .X(_01390_));
 nand2_1 _21156_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[15] ),
    .B(_03402_),
    .Y(_05832_));
 or2_1 _21157_ (.A(\digitop_pav2.aes128_inst.aes128_regs.key6_r[15] ),
    .B(_03402_),
    .X(_05833_));
 a311o_1 _21158_ (.A1(net442),
    .A2(_05832_),
    .A3(_05833_),
    .B1(net358),
    .C1(net343),
    .X(_05834_));
 o22a_1 _21159_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key6_r[15] ),
    .A2(net309),
    .B1(_05834_),
    .B2(_05507_),
    .X(_01391_));
 nor2_1 _21160_ (.A(_11214_),
    .B(net344),
    .Y(_05835_));
 o21ai_1 _21161_ (.A1(net408),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[0] ),
    .B1(net305),
    .Y(_05836_));
 a31o_1 _21162_ (.A1(net454),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[0] ),
    .A3(_07219_),
    .B1(_05442_),
    .X(_05837_));
 a22o_1 _21163_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[0] ),
    .A2(_05836_),
    .B1(_05837_),
    .B2(net305),
    .X(_01392_));
 o21ai_1 _21164_ (.A1(net407),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[1] ),
    .B1(net305),
    .Y(_05838_));
 a31o_1 _21165_ (.A1(net453),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[1] ),
    .A3(_07220_),
    .B1(_05446_),
    .X(_05839_));
 a22o_1 _21166_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[1] ),
    .A2(_05838_),
    .B1(_05839_),
    .B2(net305),
    .X(_01393_));
 o21ai_1 _21167_ (.A1(net407),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[2] ),
    .B1(net305),
    .Y(_05840_));
 a31o_1 _21168_ (.A1(net450),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[2] ),
    .A3(_07221_),
    .B1(_05451_),
    .X(_05841_));
 a22o_1 _21169_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[2] ),
    .A2(_05840_),
    .B1(_05841_),
    .B2(net305),
    .X(_01394_));
 o21ai_1 _21170_ (.A1(net409),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[3] ),
    .B1(net307),
    .Y(_05842_));
 a31o_1 _21171_ (.A1(net455),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[3] ),
    .A3(_07222_),
    .B1(_05456_),
    .X(_05843_));
 a22o_1 _21172_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[3] ),
    .A2(_05842_),
    .B1(_05843_),
    .B2(net307),
    .X(_01395_));
 o21ai_1 _21173_ (.A1(net409),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[4] ),
    .B1(net305),
    .Y(_05844_));
 a31o_1 _21174_ (.A1(net456),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[4] ),
    .A3(_07223_),
    .B1(_05460_),
    .X(_05845_));
 a22o_1 _21175_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[4] ),
    .A2(_05844_),
    .B1(_05845_),
    .B2(net307),
    .X(_01396_));
 o21ai_1 _21176_ (.A1(net409),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[5] ),
    .B1(net307),
    .Y(_05846_));
 a31o_1 _21177_ (.A1(net457),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[5] ),
    .A3(_07224_),
    .B1(_05465_),
    .X(_05847_));
 a22o_1 _21178_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[5] ),
    .A2(_05846_),
    .B1(_05847_),
    .B2(net305),
    .X(_01397_));
 o21ai_1 _21179_ (.A1(net408),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[6] ),
    .B1(net305),
    .Y(_05848_));
 a31o_1 _21180_ (.A1(net452),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[6] ),
    .A3(_07225_),
    .B1(_05470_),
    .X(_05849_));
 a22o_1 _21181_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[6] ),
    .A2(_05848_),
    .B1(_05849_),
    .B2(net305),
    .X(_01398_));
 o21ai_1 _21182_ (.A1(net405),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[7] ),
    .B1(net306),
    .Y(_05850_));
 a31o_1 _21183_ (.A1(net446),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[7] ),
    .A3(_07226_),
    .B1(_05473_),
    .X(_05851_));
 a22o_1 _21184_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[7] ),
    .A2(_05850_),
    .B1(_05851_),
    .B2(net306),
    .X(_01399_));
 o21ai_1 _21185_ (.A1(net411),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[8] ),
    .B1(net308),
    .Y(_05852_));
 a31o_1 _21186_ (.A1(net463),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[8] ),
    .A3(_07211_),
    .B1(_05477_),
    .X(_05853_));
 a22o_1 _21187_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[8] ),
    .A2(_05852_),
    .B1(_05853_),
    .B2(net308),
    .X(_01400_));
 o21ai_1 _21188_ (.A1(net405),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[9] ),
    .B1(net306),
    .Y(_05854_));
 a31o_1 _21189_ (.A1(net442),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[9] ),
    .A3(_07212_),
    .B1(_05480_),
    .X(_05855_));
 a22o_1 _21190_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[9] ),
    .A2(_05854_),
    .B1(_05855_),
    .B2(net306),
    .X(_01401_));
 o21ai_1 _21191_ (.A1(net406),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[10] ),
    .B1(net306),
    .Y(_05856_));
 a31o_1 _21192_ (.A1(net448),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[10] ),
    .A3(_07213_),
    .B1(_05484_),
    .X(_05857_));
 a22o_1 _21193_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[10] ),
    .A2(_05856_),
    .B1(_05857_),
    .B2(net306),
    .X(_01402_));
 o21ai_1 _21194_ (.A1(net411),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[11] ),
    .B1(net308),
    .Y(_05858_));
 a31o_1 _21195_ (.A1(net463),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[11] ),
    .A3(_07214_),
    .B1(_05489_),
    .X(_05859_));
 a22o_1 _21196_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[11] ),
    .A2(_05858_),
    .B1(_05859_),
    .B2(net308),
    .X(_01403_));
 o21ai_1 _21197_ (.A1(net411),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[12] ),
    .B1(net308),
    .Y(_05860_));
 a31o_1 _21198_ (.A1(net463),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[12] ),
    .A3(_07215_),
    .B1(_05494_),
    .X(_05861_));
 a22o_1 _21199_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[12] ),
    .A2(_05860_),
    .B1(_05861_),
    .B2(net308),
    .X(_01404_));
 o21ai_1 _21200_ (.A1(net410),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[13] ),
    .B1(net308),
    .Y(_05862_));
 a31o_1 _21201_ (.A1(net463),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[13] ),
    .A3(_07216_),
    .B1(_05499_),
    .X(_05863_));
 a22o_1 _21202_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[13] ),
    .A2(_05862_),
    .B1(_05863_),
    .B2(net308),
    .X(_01405_));
 o21ai_1 _21203_ (.A1(net406),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[14] ),
    .B1(net306),
    .Y(_05864_));
 a31o_1 _21204_ (.A1(net448),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[14] ),
    .A3(_07217_),
    .B1(_05504_),
    .X(_05865_));
 a22o_1 _21205_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[14] ),
    .A2(_05864_),
    .B1(_05865_),
    .B2(net306),
    .X(_01406_));
 o21ai_1 _21206_ (.A1(net406),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[15] ),
    .B1(net306),
    .Y(_05866_));
 a31o_1 _21207_ (.A1(net448),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[15] ),
    .A3(_07218_),
    .B1(_05507_),
    .X(_05867_));
 a22o_1 _21208_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.key5_r[15] ),
    .A2(_05866_),
    .B1(_05867_),
    .B2(net306),
    .X(_01407_));
 and3_4 _21209_ (.A(_11197_),
    .B(_03619_),
    .C(_05531_),
    .X(_05868_));
 nand3_4 _21210_ (.A(_11197_),
    .B(_03619_),
    .C(_05531_),
    .Y(_05869_));
 xor2_1 _21211_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[0] ),
    .X(_05870_));
 o21ai_1 _21212_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[0] ),
    .B1(net433),
    .Y(_05871_));
 a21oi_1 _21213_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[0] ),
    .B1(_05871_),
    .Y(_05872_));
 a211o_1 _21214_ (.A1(net419),
    .A2(_05870_),
    .B1(_05872_),
    .C1(_05869_),
    .X(_05873_));
 o32a_1 _21215_ (.A1(_11393_),
    .A2(_11476_),
    .A3(_05873_),
    .B1(_05868_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[0] ),
    .X(_01408_));
 o21ai_1 _21216_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[1] ),
    .B1(net432),
    .Y(_05874_));
 a21oi_1 _21217_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[1] ),
    .B1(_05874_),
    .Y(_05875_));
 or2_1 _21218_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[1] ),
    .X(_05876_));
 nand2_1 _21219_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[1] ),
    .Y(_05877_));
 a31o_1 _21220_ (.A1(net418),
    .A2(_05876_),
    .A3(_05877_),
    .B1(_05875_),
    .X(_05878_));
 or4_1 _21221_ (.A(_02182_),
    .B(_02224_),
    .C(_05869_),
    .D(_05878_),
    .X(_05879_));
 o22a_1 _21222_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[1] ),
    .A2(_05868_),
    .B1(_05879_),
    .B2(_02192_),
    .X(_01409_));
 o21ai_1 _21223_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[2] ),
    .B1(net435),
    .Y(_05880_));
 a21oi_1 _21224_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[2] ),
    .B1(_05880_),
    .Y(_05881_));
 xor2_1 _21225_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[2] ),
    .X(_05882_));
 a211o_1 _21226_ (.A1(net421),
    .A2(_05882_),
    .B1(_05881_),
    .C1(_05869_),
    .X(_05883_));
 o32a_1 _21227_ (.A1(_02265_),
    .A2(_02305_),
    .A3(_05883_),
    .B1(_05868_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ),
    .X(_01410_));
 o21ai_1 _21228_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[3] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[3] ),
    .B1(net436),
    .Y(_05884_));
 a21oi_1 _21229_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[3] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[3] ),
    .B1(_05884_),
    .Y(_05885_));
 or2_1 _21230_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[3] ),
    .X(_05886_));
 nand2_1 _21231_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[3] ),
    .Y(_05887_));
 a31o_1 _21232_ (.A1(net422),
    .A2(_05886_),
    .A3(_05887_),
    .B1(_05885_),
    .X(_05888_));
 or4_1 _21233_ (.A(_02339_),
    .B(_02382_),
    .C(_05869_),
    .D(_05888_),
    .X(_05889_));
 o22a_1 _21234_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[3] ),
    .A2(_05868_),
    .B1(_05889_),
    .B2(_02354_),
    .X(_01411_));
 or2_1 _21235_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[4] ),
    .X(_05890_));
 nand2_1 _21236_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[4] ),
    .Y(_05891_));
 o21ai_1 _21237_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[4] ),
    .B1(net440),
    .Y(_05892_));
 a21oi_1 _21238_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[4] ),
    .B1(_05892_),
    .Y(_05893_));
 a31o_1 _21239_ (.A1(net424),
    .A2(_05890_),
    .A3(_05891_),
    .B1(_05893_),
    .X(_05894_));
 or4_1 _21240_ (.A(_02413_),
    .B(_02451_),
    .C(_05869_),
    .D(_05894_),
    .X(_05895_));
 o22a_1 _21241_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[4] ),
    .A2(_05868_),
    .B1(_05895_),
    .B2(_02423_),
    .X(_01412_));
 o21ai_1 _21242_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[5] ),
    .B1(net437),
    .Y(_05896_));
 a21oi_1 _21243_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[5] ),
    .B1(_05896_),
    .Y(_05897_));
 or2_1 _21244_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[5] ),
    .X(_05898_));
 nand2_1 _21245_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[5] ),
    .Y(_05899_));
 a31o_1 _21246_ (.A1(net423),
    .A2(_05898_),
    .A3(_05899_),
    .B1(_05897_),
    .X(_05900_));
 or4_1 _21247_ (.A(_02482_),
    .B(_02522_),
    .C(_05869_),
    .D(_05900_),
    .X(_05901_));
 o22a_1 _21248_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[5] ),
    .A2(_05868_),
    .B1(_05901_),
    .B2(_02511_),
    .X(_01413_));
 or2_1 _21249_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[6] ),
    .X(_05902_));
 nand2_1 _21250_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[6] ),
    .Y(_05903_));
 or2_1 _21251_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[6] ),
    .X(_05904_));
 nand2_1 _21252_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[6] ),
    .Y(_05905_));
 a311o_1 _21253_ (.A1(net433),
    .A2(_05904_),
    .A3(_05905_),
    .B1(_02562_),
    .C1(_05869_),
    .X(_05906_));
 a31o_1 _21254_ (.A1(net421),
    .A2(_05902_),
    .A3(_05903_),
    .B1(_05906_),
    .X(_05907_));
 o32a_1 _21255_ (.A1(_02552_),
    .A2(_02590_),
    .A3(_05907_),
    .B1(_05868_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state0_r[6] ),
    .X(_01414_));
 o21ai_1 _21256_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[7] ),
    .B1(net430),
    .Y(_05908_));
 a21oi_1 _21257_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key0_r[7] ),
    .B1(_05908_),
    .Y(_05909_));
 or2_1 _21258_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[7] ),
    .X(_05910_));
 nand2_1 _21259_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key0_r[7] ),
    .Y(_05911_));
 a31o_1 _21260_ (.A1(net415),
    .A2(_05910_),
    .A3(_05911_),
    .B1(_05909_),
    .X(_05912_));
 or4_1 _21261_ (.A(_02616_),
    .B(_02651_),
    .C(_05869_),
    .D(_05912_),
    .X(_05913_));
 o22a_1 _21262_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ),
    .A2(_05868_),
    .B1(_05913_),
    .B2(_02626_),
    .X(_01415_));
 and3_1 _21263_ (.A(_11198_),
    .B(_03425_),
    .C(_03578_),
    .X(_05914_));
 and2_2 _21264_ (.A(_03579_),
    .B(_05914_),
    .X(_05915_));
 nand2_2 _21265_ (.A(_03579_),
    .B(_05914_),
    .Y(_05916_));
 nand2_1 _21266_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[8] ),
    .Y(_05917_));
 or2_1 _21267_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[8] ),
    .X(_05918_));
 a311o_1 _21268_ (.A1(net401),
    .A2(_05917_),
    .A3(_05918_),
    .B1(_03026_),
    .C1(_05916_),
    .X(_05919_));
 o32a_1 _21269_ (.A1(_02996_),
    .A2(_03436_),
    .A3(_05919_),
    .B1(_05915_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[8] ),
    .X(_01416_));
 o21ai_1 _21270_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[9] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[9] ),
    .B1(net401),
    .Y(_05920_));
 a21oi_1 _21271_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[9] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[9] ),
    .B1(_05920_),
    .Y(_05921_));
 or4_1 _21272_ (.A(_03082_),
    .B(_03444_),
    .C(_05916_),
    .D(_05921_),
    .X(_05922_));
 o22a_1 _21273_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[9] ),
    .A2(_05915_),
    .B1(_05922_),
    .B2(_03101_),
    .X(_01417_));
 or2_1 _21274_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[10] ),
    .X(_05923_));
 nand2_1 _21275_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[10] ),
    .Y(_05924_));
 a311o_1 _21276_ (.A1(net400),
    .A2(_05923_),
    .A3(_05924_),
    .B1(_03162_),
    .C1(_05916_),
    .X(_05925_));
 o32a_1 _21277_ (.A1(_03150_),
    .A2(_03449_),
    .A3(_05925_),
    .B1(_05915_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[10] ),
    .X(_01418_));
 o21ai_1 _21278_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[11] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[11] ),
    .B1(net402),
    .Y(_05926_));
 a21oi_1 _21279_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[11] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key1_r[11] ),
    .B1(_05926_),
    .Y(_05927_));
 or4_1 _21280_ (.A(_03202_),
    .B(_03461_),
    .C(_05916_),
    .D(_05927_),
    .X(_05928_));
 o22a_1 _21281_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[11] ),
    .A2(_05915_),
    .B1(_05928_),
    .B2(_03217_),
    .X(_01419_));
 nand2_1 _21282_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[12] ),
    .Y(_05929_));
 or2_1 _21283_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[12] ),
    .X(_05930_));
 a311o_1 _21284_ (.A1(net401),
    .A2(_05929_),
    .A3(_05930_),
    .B1(_03269_),
    .C1(_05916_),
    .X(_05931_));
 o32a_1 _21285_ (.A1(_03255_),
    .A2(_03469_),
    .A3(_05931_),
    .B1(_05915_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[12] ),
    .X(_01420_));
 nand2_1 _21286_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[13] ),
    .Y(_05932_));
 or2_1 _21287_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[13] ),
    .X(_05933_));
 a311o_1 _21288_ (.A1(net401),
    .A2(_05932_),
    .A3(_05933_),
    .B1(_03315_),
    .C1(_05916_),
    .X(_05934_));
 o32a_1 _21289_ (.A1(_03303_),
    .A2(_03477_),
    .A3(_05934_),
    .B1(_05915_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[13] ),
    .X(_01421_));
 or2_1 _21290_ (.A(_03363_),
    .B(_03482_),
    .X(_05935_));
 or2_1 _21291_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[14] ),
    .X(_05936_));
 nand2_1 _21292_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[14] ),
    .Y(_05937_));
 a31o_1 _21293_ (.A1(net399),
    .A2(_05936_),
    .A3(_05937_),
    .B1(_05916_),
    .X(_05938_));
 o22a_1 _21294_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state1_r[14] ),
    .A2(_05915_),
    .B1(_05935_),
    .B2(_05938_),
    .X(_01422_));
 or2_1 _21295_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[15] ),
    .X(_05939_));
 nand2_1 _21296_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state1_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key1_r[15] ),
    .Y(_05940_));
 a31o_1 _21297_ (.A1(net399),
    .A2(_05939_),
    .A3(_05940_),
    .B1(_05916_),
    .X(_05941_));
 o32a_1 _21298_ (.A1(_03412_),
    .A2(_03491_),
    .A3(_05941_),
    .B1(_05915_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state1_r[15] ),
    .X(_01423_));
 and3_2 _21299_ (.A(_11203_),
    .B(_02824_),
    .C(_05531_),
    .X(_05942_));
 nand3_4 _21300_ (.A(_11203_),
    .B(_02824_),
    .C(_05531_),
    .Y(_05943_));
 or2_1 _21301_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[8] ),
    .X(_05944_));
 nand2_1 _21302_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[8] ),
    .Y(_05945_));
 or2_1 _21303_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[8] ),
    .X(_05946_));
 nand2_1 _21304_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[8] ),
    .Y(_05947_));
 a311o_1 _21305_ (.A1(net416),
    .A2(_05946_),
    .A3(_05947_),
    .B1(_03026_),
    .C1(_05943_),
    .X(_05948_));
 a31o_1 _21306_ (.A1(net431),
    .A2(_05944_),
    .A3(_05945_),
    .B1(_05948_),
    .X(_05949_));
 a31o_1 _21307_ (.A1(net468),
    .A2(_03029_),
    .A3(_03030_),
    .B1(_05949_),
    .X(_05950_));
 o22a_1 _21308_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[8] ),
    .A2(_05942_),
    .B1(_05950_),
    .B2(_02996_),
    .X(_01424_));
 o21ai_1 _21309_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[9] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[9] ),
    .B1(net429),
    .Y(_05951_));
 a21oi_1 _21310_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[9] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[9] ),
    .B1(_05951_),
    .Y(_05952_));
 or2_1 _21311_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[9] ),
    .X(_05953_));
 nand2_1 _21312_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[9] ),
    .Y(_05954_));
 a31o_1 _21313_ (.A1(net414),
    .A2(_05953_),
    .A3(_05954_),
    .B1(_05952_),
    .X(_05955_));
 or4b_1 _21314_ (.A(_03082_),
    .B(_05943_),
    .C(_05955_),
    .D_N(_03106_),
    .X(_05956_));
 o22a_1 _21315_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[9] ),
    .A2(_05942_),
    .B1(_05956_),
    .B2(_03101_),
    .X(_01425_));
 or2_1 _21316_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[10] ),
    .X(_05957_));
 nand2_1 _21317_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[10] ),
    .Y(_05958_));
 or2_1 _21318_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[10] ),
    .X(_05959_));
 nand2_1 _21319_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[10] ),
    .Y(_05960_));
 a311o_1 _21320_ (.A1(net416),
    .A2(_05957_),
    .A3(_05958_),
    .B1(_03162_),
    .C1(_05943_),
    .X(_05961_));
 a31o_1 _21321_ (.A1(net431),
    .A2(_05959_),
    .A3(_05960_),
    .B1(_05961_),
    .X(_05962_));
 o32a_1 _21322_ (.A1(_03150_),
    .A2(_03171_),
    .A3(_05962_),
    .B1(_05942_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[10] ),
    .X(_01426_));
 or2_1 _21323_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[11] ),
    .X(_05963_));
 nand2_1 _21324_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[11] ),
    .Y(_05964_));
 or2_1 _21325_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[11] ),
    .X(_05965_));
 nand2_1 _21326_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[11] ),
    .Y(_05966_));
 a31o_1 _21327_ (.A1(net425),
    .A2(_05965_),
    .A3(_05966_),
    .B1(_05943_),
    .X(_05967_));
 a311o_1 _21328_ (.A1(net438),
    .A2(_05963_),
    .A3(_05964_),
    .B1(_05967_),
    .C1(_03217_),
    .X(_05968_));
 o32a_1 _21329_ (.A1(_03202_),
    .A2(_03223_),
    .A3(_05968_),
    .B1(_05942_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[11] ),
    .X(_01427_));
 or2_1 _21330_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[12] ),
    .X(_05969_));
 nand2_1 _21331_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state2_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[12] ),
    .Y(_05970_));
 or2_1 _21332_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[12] ),
    .X(_05971_));
 nand2_1 _21333_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[12] ),
    .Y(_05972_));
 a311o_1 _21334_ (.A1(net416),
    .A2(_05971_),
    .A3(_05972_),
    .B1(_03269_),
    .C1(_05943_),
    .X(_05973_));
 a31o_1 _21335_ (.A1(net438),
    .A2(_05969_),
    .A3(_05970_),
    .B1(_05973_),
    .X(_05974_));
 o32a_1 _21336_ (.A1(_03255_),
    .A2(_03274_),
    .A3(_05974_),
    .B1(_05942_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[12] ),
    .X(_01428_));
 o21ai_1 _21337_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[13] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[13] ),
    .B1(net439),
    .Y(_05975_));
 a21oi_1 _21338_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[13] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[13] ),
    .B1(_05975_),
    .Y(_05976_));
 or2_1 _21339_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[13] ),
    .X(_05977_));
 nand2_1 _21340_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[13] ),
    .Y(_05978_));
 a311o_1 _21341_ (.A1(net427),
    .A2(_05977_),
    .A3(_05978_),
    .B1(_05943_),
    .C1(_05976_),
    .X(_05979_));
 o32a_1 _21342_ (.A1(_03303_),
    .A2(_03526_),
    .A3(_05979_),
    .B1(_05942_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[13] ),
    .X(_01429_));
 o21ai_1 _21343_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[14] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[14] ),
    .B1(net429),
    .Y(_05980_));
 a21oi_1 _21344_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[14] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[14] ),
    .B1(_05980_),
    .Y(_05981_));
 or2_1 _21345_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[14] ),
    .X(_05982_));
 nand2_1 _21346_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[14] ),
    .Y(_05983_));
 a31o_1 _21347_ (.A1(net414),
    .A2(_05982_),
    .A3(_05983_),
    .B1(_05981_),
    .X(_05984_));
 or3_1 _21348_ (.A(_03363_),
    .B(_05943_),
    .C(_05984_),
    .X(_05985_));
 o32a_1 _21349_ (.A1(_03353_),
    .A2(_03374_),
    .A3(_05985_),
    .B1(_05942_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[14] ),
    .X(_01430_));
 o21ai_1 _21350_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[15] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[15] ),
    .B1(net430),
    .Y(_05986_));
 a21oi_1 _21351_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state2_r[15] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key2_r[15] ),
    .B1(_05986_),
    .Y(_05987_));
 xor2_1 _21352_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key2_r[15] ),
    .X(_05988_));
 a2111o_1 _21353_ (.A1(net415),
    .A2(_05988_),
    .B1(_05987_),
    .C1(_05943_),
    .D1(_03412_),
    .X(_05989_));
 o32a_1 _21354_ (.A1(_03403_),
    .A2(_03421_),
    .A3(_05989_),
    .B1(_05942_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state2_r[15] ),
    .X(_01431_));
 and4b_4 _21355_ (.A_N(_11194_),
    .B(_02823_),
    .C(_03425_),
    .D(_03535_),
    .X(_05990_));
 a2111o_4 _21356_ (.A1(net468),
    .A2(_11444_),
    .B1(_03424_),
    .C1(_03536_),
    .D1(_11194_),
    .X(_05991_));
 nand2_1 _21357_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[8] ),
    .Y(_05992_));
 or2_1 _21358_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[8] ),
    .X(_05993_));
 a311o_1 _21359_ (.A1(net401),
    .A2(_05992_),
    .A3(_05993_),
    .B1(_03026_),
    .C1(_05991_),
    .X(_05994_));
 o32a_1 _21360_ (.A1(_02996_),
    .A2(_03436_),
    .A3(_05994_),
    .B1(_05990_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[8] ),
    .X(_01432_));
 nand2_1 _21361_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[9] ),
    .Y(_05995_));
 or2_1 _21362_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[9] ),
    .X(_05996_));
 a311o_1 _21363_ (.A1(net401),
    .A2(_05995_),
    .A3(_05996_),
    .B1(_03101_),
    .C1(_05991_),
    .X(_05997_));
 o32a_1 _21364_ (.A1(_03082_),
    .A2(_03444_),
    .A3(_05997_),
    .B1(_05990_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[9] ),
    .X(_01433_));
 or2_1 _21365_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[10] ),
    .X(_05998_));
 nand2_1 _21366_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[10] ),
    .Y(_05999_));
 a311o_1 _21367_ (.A1(net400),
    .A2(_05998_),
    .A3(_05999_),
    .B1(_03162_),
    .C1(_05991_),
    .X(_06000_));
 o32a_1 _21368_ (.A1(_03150_),
    .A2(_03449_),
    .A3(_06000_),
    .B1(_05990_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[10] ),
    .X(_01434_));
 nand2_1 _21369_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[11] ),
    .Y(_06001_));
 or2_1 _21370_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[11] ),
    .X(_06002_));
 a311o_1 _21371_ (.A1(net401),
    .A2(_06001_),
    .A3(_06002_),
    .B1(_03217_),
    .C1(_05991_),
    .X(_06003_));
 o32a_1 _21372_ (.A1(_03202_),
    .A2(_03461_),
    .A3(_06003_),
    .B1(_05990_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[11] ),
    .X(_01435_));
 nand2_1 _21373_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[12] ),
    .Y(_06004_));
 or2_1 _21374_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[12] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[12] ),
    .X(_06005_));
 a311o_1 _21375_ (.A1(net401),
    .A2(_06004_),
    .A3(_06005_),
    .B1(_03269_),
    .C1(_05991_),
    .X(_06006_));
 o32a_1 _21376_ (.A1(_03255_),
    .A2(_03469_),
    .A3(_06006_),
    .B1(_05990_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[12] ),
    .X(_01436_));
 nand2_1 _21377_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[13] ),
    .Y(_06007_));
 or2_1 _21378_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[13] ),
    .X(_06008_));
 a311o_1 _21379_ (.A1(net401),
    .A2(_06007_),
    .A3(_06008_),
    .B1(_03315_),
    .C1(_05991_),
    .X(_06009_));
 o32a_1 _21380_ (.A1(_03303_),
    .A2(_03477_),
    .A3(_06009_),
    .B1(_05990_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state3_r[13] ),
    .X(_01437_));
 or2_1 _21381_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[14] ),
    .X(_06010_));
 nand2_1 _21382_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[14] ),
    .Y(_06011_));
 a31o_1 _21383_ (.A1(net399),
    .A2(_06010_),
    .A3(_06011_),
    .B1(_05991_),
    .X(_06012_));
 o22a_1 _21384_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[14] ),
    .A2(_05990_),
    .B1(_06012_),
    .B2(_05935_),
    .X(_01438_));
 or2_1 _21385_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[15] ),
    .X(_06013_));
 nand2_1 _21386_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state3_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key3_r[15] ),
    .Y(_06014_));
 a311o_1 _21387_ (.A1(net399),
    .A2(_06013_),
    .A3(_06014_),
    .B1(_03412_),
    .C1(_05991_),
    .X(_06015_));
 o22a_1 _21388_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state3_r[15] ),
    .A2(_05990_),
    .B1(_06015_),
    .B2(_03491_),
    .X(_01439_));
 nand2_1 _21389_ (.A(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[0] ),
    .B(_10786_),
    .Y(_06016_));
 o221a_1 _21390_ (.A1(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[0] ),
    .A2(_10751_),
    .B1(_10783_),
    .B2(_10750_),
    .C1(_06016_),
    .X(_01440_));
 a211o_1 _21391_ (.A1(_11199_),
    .A2(_11212_),
    .B1(_10744_),
    .C1(_10749_),
    .X(_06017_));
 o221ai_1 _21392_ (.A1(_07105_),
    .A2(_10751_),
    .B1(_10780_),
    .B2(_10750_),
    .C1(_06017_),
    .Y(_01441_));
 nor2_1 _21393_ (.A(_10744_),
    .B(_11210_),
    .Y(_06018_));
 xnor2_1 _21394_ (.A(_07106_),
    .B(_06018_),
    .Y(_06019_));
 mux2_1 _21395_ (.A0(_10777_),
    .A1(_06019_),
    .S(_10750_),
    .X(_01442_));
 and3_2 _21396_ (.A(net334),
    .B(_03425_),
    .C(_05531_),
    .X(_06020_));
 nand3_4 _21397_ (.A(net334),
    .B(_03425_),
    .C(_05531_),
    .Y(_06021_));
 nand2_1 _21398_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[8] ),
    .Y(_06022_));
 or2_1 _21399_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[8] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[8] ),
    .X(_06023_));
 a311o_1 _21400_ (.A1(net402),
    .A2(_06022_),
    .A3(_06023_),
    .B1(_03026_),
    .C1(_06021_),
    .X(_06024_));
 o32a_1 _21401_ (.A1(_02996_),
    .A2(_03436_),
    .A3(_06024_),
    .B1(_06020_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[8] ),
    .X(_01443_));
 nand2_1 _21402_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[9] ),
    .Y(_06025_));
 or2_1 _21403_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[9] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[9] ),
    .X(_06026_));
 a311o_1 _21404_ (.A1(net399),
    .A2(_06025_),
    .A3(_06026_),
    .B1(_03101_),
    .C1(_06021_),
    .X(_06027_));
 o32a_1 _21405_ (.A1(_03082_),
    .A2(_03444_),
    .A3(_06027_),
    .B1(_06020_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[9] ),
    .X(_01444_));
 nand2_1 _21406_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[10] ),
    .Y(_06028_));
 or2_1 _21407_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[10] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[10] ),
    .X(_06029_));
 a311o_1 _21408_ (.A1(net399),
    .A2(_06028_),
    .A3(_06029_),
    .B1(_03162_),
    .C1(_06021_),
    .X(_06030_));
 o32a_1 _21409_ (.A1(_03150_),
    .A2(_03449_),
    .A3(_06030_),
    .B1(_06020_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[10] ),
    .X(_01445_));
 nand2_1 _21410_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[11] ),
    .Y(_06031_));
 or2_1 _21411_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[11] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[11] ),
    .X(_06032_));
 a311o_1 _21412_ (.A1(net402),
    .A2(_06031_),
    .A3(_06032_),
    .B1(_03217_),
    .C1(_06021_),
    .X(_06033_));
 o32a_1 _21413_ (.A1(_03202_),
    .A2(_03461_),
    .A3(_06033_),
    .B1(_06020_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[11] ),
    .X(_01446_));
 o21ai_1 _21414_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[12] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[12] ),
    .B1(_11222_),
    .Y(_06034_));
 a21oi_1 _21415_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[12] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key7_r[12] ),
    .B1(_06034_),
    .Y(_06035_));
 or4_1 _21416_ (.A(_03255_),
    .B(_03469_),
    .C(_06021_),
    .D(_06035_),
    .X(_06036_));
 o22a_1 _21417_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[12] ),
    .A2(_06020_),
    .B1(_06036_),
    .B2(_03269_),
    .X(_01447_));
 nand2_1 _21418_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[13] ),
    .Y(_06037_));
 or2_1 _21419_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[13] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[13] ),
    .X(_06038_));
 a311o_1 _21420_ (.A1(net402),
    .A2(_06037_),
    .A3(_06038_),
    .B1(_03315_),
    .C1(_06021_),
    .X(_06039_));
 o32a_1 _21421_ (.A1(_03303_),
    .A2(_03477_),
    .A3(_06039_),
    .B1(_06020_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[13] ),
    .X(_01448_));
 or2_1 _21422_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[14] ),
    .X(_06040_));
 nand2_1 _21423_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[14] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[14] ),
    .Y(_06041_));
 a31o_1 _21424_ (.A1(net400),
    .A2(_06040_),
    .A3(_06041_),
    .B1(_06021_),
    .X(_06042_));
 o22a_1 _21425_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state7_r[14] ),
    .A2(_06020_),
    .B1(_06042_),
    .B2(_05935_),
    .X(_01449_));
 or2_1 _21426_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[15] ),
    .X(_06043_));
 nand2_1 _21427_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state7_r[15] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key7_r[15] ),
    .Y(_06044_));
 a31o_1 _21428_ (.A1(net399),
    .A2(_06043_),
    .A3(_06044_),
    .B1(_06021_),
    .X(_06045_));
 o32a_1 _21429_ (.A1(_03412_),
    .A2(_03491_),
    .A3(_06045_),
    .B1(_06020_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state7_r[15] ),
    .X(_01450_));
 and3_4 _21430_ (.A(_11197_),
    .B(_02822_),
    .C(_03422_),
    .X(_06046_));
 nand3_4 _21431_ (.A(_11197_),
    .B(_02822_),
    .C(_03422_),
    .Y(_06047_));
 o21ai_1 _21432_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[0] ),
    .B1(net433),
    .Y(_06048_));
 a21oi_1 _21433_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[0] ),
    .B1(_06048_),
    .Y(_06049_));
 or2_1 _21434_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[0] ),
    .X(_06050_));
 nand2_1 _21435_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[0] ),
    .Y(_06051_));
 a311o_1 _21436_ (.A1(net419),
    .A2(_06050_),
    .A3(_06051_),
    .B1(_06047_),
    .C1(_06049_),
    .X(_06052_));
 o32a_1 _21437_ (.A1(_11393_),
    .A2(_11476_),
    .A3(_06052_),
    .B1(_06046_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[0] ),
    .X(_01451_));
 or2_1 _21438_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[1] ),
    .X(_06053_));
 nand2_1 _21439_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[1] ),
    .Y(_06054_));
 o21ai_1 _21440_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[1] ),
    .B1(net432),
    .Y(_06055_));
 a21oi_1 _21441_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[1] ),
    .B1(_06055_),
    .Y(_06056_));
 a31o_1 _21442_ (.A1(net418),
    .A2(_06053_),
    .A3(_06054_),
    .B1(_06056_),
    .X(_06057_));
 or4_1 _21443_ (.A(_02182_),
    .B(_02224_),
    .C(_06047_),
    .D(_06057_),
    .X(_06058_));
 o22a_1 _21444_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[1] ),
    .A2(_06046_),
    .B1(_06058_),
    .B2(_02192_),
    .X(_01452_));
 o21ai_1 _21445_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[2] ),
    .B1(net435),
    .Y(_06059_));
 a21oi_1 _21446_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[2] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[2] ),
    .B1(_06059_),
    .Y(_06060_));
 or2_1 _21447_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[2] ),
    .X(_06061_));
 nand2_1 _21448_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[2] ),
    .Y(_06062_));
 a311o_1 _21449_ (.A1(net421),
    .A2(_06061_),
    .A3(_06062_),
    .B1(_06047_),
    .C1(_06060_),
    .X(_06063_));
 o32a_1 _21450_ (.A1(_02265_),
    .A2(_02305_),
    .A3(_06063_),
    .B1(_06046_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[2] ),
    .X(_01453_));
 o21ai_1 _21451_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[3] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[3] ),
    .B1(net436),
    .Y(_06064_));
 a21oi_1 _21452_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[3] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[3] ),
    .B1(_06064_),
    .Y(_06065_));
 or2_1 _21453_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[3] ),
    .X(_06066_));
 nand2_1 _21454_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[3] ),
    .Y(_06067_));
 a31o_1 _21455_ (.A1(net422),
    .A2(_06066_),
    .A3(_06067_),
    .B1(_06065_),
    .X(_06068_));
 or4_1 _21456_ (.A(_02339_),
    .B(_02382_),
    .C(_06047_),
    .D(_06068_),
    .X(_06069_));
 o22a_1 _21457_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[3] ),
    .A2(_06046_),
    .B1(_06069_),
    .B2(_02354_),
    .X(_01454_));
 or2_1 _21458_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[4] ),
    .X(_06070_));
 nand2_1 _21459_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[4] ),
    .Y(_06071_));
 o21ai_1 _21460_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[4] ),
    .B1(net437),
    .Y(_06072_));
 a21oi_1 _21461_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[4] ),
    .B1(_06072_),
    .Y(_06073_));
 a31o_1 _21462_ (.A1(net423),
    .A2(_06070_),
    .A3(_06071_),
    .B1(_06073_),
    .X(_06074_));
 or4_1 _21463_ (.A(_02413_),
    .B(_02451_),
    .C(_06047_),
    .D(_06074_),
    .X(_06075_));
 o22a_1 _21464_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[4] ),
    .A2(_06046_),
    .B1(_06075_),
    .B2(_02423_),
    .X(_01455_));
 o21ai_1 _21465_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[5] ),
    .B1(net437),
    .Y(_06076_));
 a21oi_1 _21466_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[5] ),
    .B1(_06076_),
    .Y(_06077_));
 or2_1 _21467_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[5] ),
    .X(_06078_));
 nand2_1 _21468_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[5] ),
    .Y(_06079_));
 a31o_1 _21469_ (.A1(net422),
    .A2(_06078_),
    .A3(_06079_),
    .B1(_06077_),
    .X(_06080_));
 or4_1 _21470_ (.A(_02482_),
    .B(_02522_),
    .C(_06047_),
    .D(_06080_),
    .X(_06081_));
 o22a_1 _21471_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[5] ),
    .A2(_06046_),
    .B1(_06081_),
    .B2(_02511_),
    .X(_01456_));
 or2_1 _21472_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[6] ),
    .X(_06082_));
 nand2_1 _21473_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[6] ),
    .Y(_06083_));
 or2_1 _21474_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[6] ),
    .X(_06084_));
 nand2_1 _21475_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[6] ),
    .Y(_06085_));
 a311o_1 _21476_ (.A1(net419),
    .A2(_06082_),
    .A3(_06083_),
    .B1(_02562_),
    .C1(_06047_),
    .X(_06086_));
 a31o_1 _21477_ (.A1(net433),
    .A2(_06084_),
    .A3(_06085_),
    .B1(_06086_),
    .X(_06087_));
 o32a_1 _21478_ (.A1(_02552_),
    .A2(_02590_),
    .A3(_06087_),
    .B1(_06046_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state6_r[6] ),
    .X(_01457_));
 o21ai_1 _21479_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[7] ),
    .B1(net430),
    .Y(_06088_));
 a21oi_1 _21480_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key6_r[7] ),
    .B1(_06088_),
    .Y(_06089_));
 or2_1 _21481_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[7] ),
    .X(_06090_));
 nand2_1 _21482_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key6_r[7] ),
    .Y(_06091_));
 a31o_1 _21483_ (.A1(net415),
    .A2(_06090_),
    .A3(_06091_),
    .B1(_06089_),
    .X(_06092_));
 or4_1 _21484_ (.A(_02616_),
    .B(_02651_),
    .C(_06047_),
    .D(_06092_),
    .X(_06093_));
 o22a_1 _21485_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[7] ),
    .A2(_06046_),
    .B1(_06093_),
    .B2(_02626_),
    .X(_01458_));
 and3_4 _21486_ (.A(_11197_),
    .B(_02823_),
    .C(_03495_),
    .X(_06094_));
 nand3_4 _21487_ (.A(_11197_),
    .B(_02823_),
    .C(_03495_),
    .Y(_06095_));
 o21ai_1 _21488_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[0] ),
    .B1(net433),
    .Y(_06096_));
 a21oi_1 _21489_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[0] ),
    .B1(_06096_),
    .Y(_06097_));
 xor2_1 _21490_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[0] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[0] ),
    .X(_06098_));
 a211o_1 _21491_ (.A1(net420),
    .A2(_06098_),
    .B1(_06097_),
    .C1(_06095_),
    .X(_06099_));
 o32a_1 _21492_ (.A1(_11393_),
    .A2(_11476_),
    .A3(_06099_),
    .B1(_06094_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ),
    .X(_01459_));
 o21ai_1 _21493_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[1] ),
    .B1(net432),
    .Y(_06100_));
 a21oi_1 _21494_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[1] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[1] ),
    .B1(_06100_),
    .Y(_06101_));
 or2_1 _21495_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[1] ),
    .X(_06102_));
 nand2_1 _21496_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[1] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[1] ),
    .Y(_06103_));
 a31o_1 _21497_ (.A1(net418),
    .A2(_06102_),
    .A3(_06103_),
    .B1(_06101_),
    .X(_06104_));
 or4_1 _21498_ (.A(_02182_),
    .B(_02224_),
    .C(_06095_),
    .D(_06104_),
    .X(_06105_));
 o22a_1 _21499_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[1] ),
    .A2(_06094_),
    .B1(_06105_),
    .B2(_02192_),
    .X(_01460_));
 or2_1 _21500_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[2] ),
    .X(_06106_));
 nand2_1 _21501_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[2] ),
    .Y(_06107_));
 or2_1 _21502_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[2] ),
    .X(_06108_));
 nand2_1 _21503_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[2] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[2] ),
    .Y(_06109_));
 a311o_1 _21504_ (.A1(net421),
    .A2(_06106_),
    .A3(_06107_),
    .B1(_02280_),
    .C1(_06095_),
    .X(_06110_));
 a31o_1 _21505_ (.A1(net435),
    .A2(_06108_),
    .A3(_06109_),
    .B1(_06110_),
    .X(_06111_));
 o32a_1 _21506_ (.A1(_02265_),
    .A2(_02304_),
    .A3(_06111_),
    .B1(_06094_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[2] ),
    .X(_01461_));
 o21ai_1 _21507_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[3] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[3] ),
    .B1(net422),
    .Y(_06112_));
 a21oi_1 _21508_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[3] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[3] ),
    .B1(_06112_),
    .Y(_06113_));
 or2_1 _21509_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[3] ),
    .X(_06114_));
 nand2_1 _21510_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[3] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[3] ),
    .Y(_06115_));
 a31o_1 _21511_ (.A1(net436),
    .A2(_06114_),
    .A3(_06115_),
    .B1(_06113_),
    .X(_06116_));
 or4_1 _21512_ (.A(_02339_),
    .B(_02382_),
    .C(_06095_),
    .D(_06116_),
    .X(_06117_));
 o22a_1 _21513_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[3] ),
    .A2(_06094_),
    .B1(_06117_),
    .B2(_02354_),
    .X(_01462_));
 o21ai_1 _21514_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[4] ),
    .B1(net437),
    .Y(_06118_));
 a21oi_1 _21515_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[4] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[4] ),
    .B1(_06118_),
    .Y(_06119_));
 or2_1 _21516_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[4] ),
    .X(_06120_));
 nand2_1 _21517_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[4] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[4] ),
    .Y(_06121_));
 a31o_1 _21518_ (.A1(net423),
    .A2(_06120_),
    .A3(_06121_),
    .B1(_06119_),
    .X(_06122_));
 or4_1 _21519_ (.A(_02413_),
    .B(_02451_),
    .C(_06095_),
    .D(_06122_),
    .X(_06123_));
 o22a_1 _21520_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[4] ),
    .A2(_06094_),
    .B1(_06123_),
    .B2(_02423_),
    .X(_01463_));
 o21ai_1 _21521_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[5] ),
    .B1(net440),
    .Y(_06124_));
 a21oi_1 _21522_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[5] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[5] ),
    .B1(_06124_),
    .Y(_06125_));
 or2_1 _21523_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[5] ),
    .X(_06126_));
 nand2_1 _21524_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[5] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[5] ),
    .Y(_06127_));
 a31o_1 _21525_ (.A1(net423),
    .A2(_06126_),
    .A3(_06127_),
    .B1(_06125_),
    .X(_06128_));
 or4_1 _21526_ (.A(_02482_),
    .B(_02522_),
    .C(_06095_),
    .D(_06128_),
    .X(_06129_));
 o22a_1 _21527_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[5] ),
    .A2(_06094_),
    .B1(_06129_),
    .B2(_02511_),
    .X(_01464_));
 xor2_1 _21528_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state6_r[6] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[6] ),
    .X(_06130_));
 o21ai_1 _21529_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[6] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[6] ),
    .B1(net433),
    .Y(_06131_));
 a21oi_1 _21530_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[6] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[6] ),
    .B1(_06131_),
    .Y(_06132_));
 a2111o_1 _21531_ (.A1(net419),
    .A2(_06130_),
    .B1(_06132_),
    .C1(_02562_),
    .D1(_06095_),
    .X(_06133_));
 o32a_1 _21532_ (.A1(_02552_),
    .A2(_02590_),
    .A3(_06133_),
    .B1(_06094_),
    .B2(\digitop_pav2.aes128_inst.aes128_regs.state4_r[6] ),
    .X(_01465_));
 o21ai_1 _21533_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[7] ),
    .B1(net415),
    .Y(_06134_));
 a21oi_1 _21534_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state6_r[7] ),
    .A2(\digitop_pav2.aes128_inst.aes128_regs.key4_r[7] ),
    .B1(_06134_),
    .Y(_06135_));
 or2_1 _21535_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[7] ),
    .X(_06136_));
 nand2_1 _21536_ (.A(\digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ),
    .B(\digitop_pav2.aes128_inst.aes128_regs.key4_r[7] ),
    .Y(_06137_));
 a31o_1 _21537_ (.A1(net430),
    .A2(_06136_),
    .A3(_06137_),
    .B1(_06135_),
    .X(_06138_));
 or4_1 _21538_ (.A(_02616_),
    .B(_02651_),
    .C(_06095_),
    .D(_06138_),
    .X(_06139_));
 o22a_1 _21539_ (.A1(\digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ),
    .A2(_06094_),
    .B1(_06139_),
    .B2(_02626_),
    .X(_01466_));
 mux2_1 _21540_ (.A0(\digitop_pav2.ack_inst.rcnt_ff[0] ),
    .A1(_07905_),
    .S(_10447_),
    .X(_01467_));
 a21o_1 _21541_ (.A1(\digitop_pav2.ack_inst.rcnt_ff[0] ),
    .A2(_10447_),
    .B1(\digitop_pav2.ack_inst.rcnt_ff[1] ),
    .X(_01468_));
 mux2_1 _21542_ (.A0(\digitop_pav2.pie_inst.fsm.pivot[0] ),
    .A1(\digitop_pav2.pie_inst.fsm.dif_pos_fix[1] ),
    .S(net475),
    .X(_01469_));
 mux2_1 _21543_ (.A0(\digitop_pav2.pie_inst.fsm.pivot[1] ),
    .A1(\digitop_pav2.pie_inst.fsm.dif_pos_fix[2] ),
    .S(net475),
    .X(_01470_));
 mux2_1 _21544_ (.A0(\digitop_pav2.pie_inst.fsm.pivot[2] ),
    .A1(\digitop_pav2.pie_inst.fsm.dif_pos_fix[3] ),
    .S(_00991_),
    .X(_01471_));
 mux2_1 _21545_ (.A0(\digitop_pav2.pie_inst.fsm.pivot[3] ),
    .A1(\digitop_pav2.pie_inst.fsm.dif_pos_fix[4] ),
    .S(net475),
    .X(_01472_));
 mux2_1 _21546_ (.A0(\digitop_pav2.pie_inst.fsm.pivot[4] ),
    .A1(\digitop_pav2.pie_inst.fsm.dif_pos_fix[5] ),
    .S(net475),
    .X(_01473_));
 mux2_1 _21547_ (.A0(\digitop_pav2.pie_inst.fsm.pivot[5] ),
    .A1(\digitop_pav2.pie_inst.fsm.dif_pos_fix[6] ),
    .S(net475),
    .X(_01474_));
 mux2_1 _21548_ (.A0(net1300),
    .A1(\digitop_pav2.pie_inst.fsm.dif_pos_fix[7] ),
    .S(net475),
    .X(_01475_));
 mux2_1 _21549_ (.A0(\digitop_pav2.pie_inst.fsm.pivot[7] ),
    .A1(\digitop_pav2.pie_inst.fsm.dif_pos_fix[8] ),
    .S(net475),
    .X(_01476_));
 mux2_1 _21550_ (.A0(\digitop_pav2.pie_inst.fsm.pivot[8] ),
    .A1(\digitop_pav2.pie_inst.fsm.dif_pos_fix[9] ),
    .S(net475),
    .X(_01477_));
 a211oi_2 _21551_ (.A1(\digitop_pav2.ack_inst.state_ff[1] ),
    .A2(_08511_),
    .B1(_07862_),
    .C1(net1234),
    .Y(_06140_));
 xnor2_1 _21552_ (.A(_07054_),
    .B(_06140_),
    .Y(_01478_));
 and3_1 _21553_ (.A(\digitop_pav2.ack_inst.cnt_ff[0] ),
    .B(net1182),
    .C(_06140_),
    .X(_06141_));
 a21oi_1 _21554_ (.A1(\digitop_pav2.ack_inst.cnt_ff[0] ),
    .A2(_06140_),
    .B1(net1182),
    .Y(_06142_));
 nor2_1 _21555_ (.A(_06141_),
    .B(_06142_),
    .Y(_01479_));
 and2_1 _21556_ (.A(\digitop_pav2.ack_inst.cnt_ff[2] ),
    .B(_06141_),
    .X(_06143_));
 xnor2_1 _21557_ (.A(_07088_),
    .B(_06141_),
    .Y(_01480_));
 xnor2_1 _21558_ (.A(_07089_),
    .B(_06143_),
    .Y(_01481_));
 mux2_1 _21559_ (.A0(net1640),
    .A1(net1082),
    .S(_02732_),
    .X(_01482_));
 mux2_1 _21560_ (.A0(net1082),
    .A1(net1080),
    .S(_02732_),
    .X(_01483_));
 mux2_1 _21561_ (.A0(net1080),
    .A1(net1078),
    .S(_02732_),
    .X(_01484_));
 mux2_1 _21562_ (.A0(net1078),
    .A1(net1076),
    .S(_02732_),
    .X(_01485_));
 mux2_1 _21563_ (.A0(net1076),
    .A1(\digitop_pav2.access_inst.access_check0.wordptr_i[4] ),
    .S(_02732_),
    .X(_01486_));
 mux2_1 _21564_ (.A0(net1074),
    .A1(net1073),
    .S(_02732_),
    .X(_01487_));
 mux2_1 _21565_ (.A0(net1073),
    .A1(net1072),
    .S(_02732_),
    .X(_01488_));
 and2_1 _21566_ (.A(_07864_),
    .B(_10447_),
    .X(_06144_));
 inv_2 _21567_ (.A(net1161),
    .Y(_06145_));
 mux2_1 _21568_ (.A0(\digitop_pav2.ack_inst.buffer_ff[0] ),
    .A1(net1135),
    .S(net1160),
    .X(_01489_));
 mux2_1 _21569_ (.A0(\digitop_pav2.ack_inst.buffer_ff[1] ),
    .A1(net1133),
    .S(net1160),
    .X(_01490_));
 mux2_1 _21570_ (.A0(\digitop_pav2.ack_inst.buffer_ff[2] ),
    .A1(net1129),
    .S(net1160),
    .X(_01491_));
 nand2_1 _21571_ (.A(_07888_),
    .B(_07905_),
    .Y(_06146_));
 a32o_1 _21572_ (.A1(net1125),
    .A2(_10447_),
    .A3(_06146_),
    .B1(_06145_),
    .B2(\digitop_pav2.ack_inst.buffer_ff[3] ),
    .X(_01492_));
 mux2_1 _21573_ (.A0(\digitop_pav2.ack_inst.buffer_ff[4] ),
    .A1(net1122),
    .S(net1160),
    .X(_01493_));
 mux2_1 _21574_ (.A0(\digitop_pav2.ack_inst.buffer_ff[5] ),
    .A1(net1119),
    .S(net1160),
    .X(_01494_));
 mux2_1 _21575_ (.A0(\digitop_pav2.ack_inst.buffer_ff[6] ),
    .A1(net1116),
    .S(net1161),
    .X(_01495_));
 mux2_1 _21576_ (.A0(\digitop_pav2.ack_inst.buffer_ff[7] ),
    .A1(net1113),
    .S(net1160),
    .X(_01496_));
 mux2_1 _21577_ (.A0(\digitop_pav2.ack_inst.buffer_ff[8] ),
    .A1(net1109),
    .S(net1161),
    .X(_01497_));
 mux2_1 _21578_ (.A0(\digitop_pav2.ack_inst.buffer_ff[9] ),
    .A1(net1105),
    .S(net1160),
    .X(_01498_));
 mux2_1 _21579_ (.A0(\digitop_pav2.ack_inst.buffer_ff[10] ),
    .A1(net1101),
    .S(net1160),
    .X(_01499_));
 mux2_1 _21580_ (.A0(\digitop_pav2.ack_inst.buffer_ff[11] ),
    .A1(net1097),
    .S(net1160),
    .X(_01500_));
 mux2_1 _21581_ (.A0(\digitop_pav2.ack_inst.buffer_ff[12] ),
    .A1(net1095),
    .S(net1161),
    .X(_01501_));
 mux2_1 _21582_ (.A0(\digitop_pav2.ack_inst.buffer_ff[13] ),
    .A1(net1092),
    .S(net1161),
    .X(_01502_));
 mux2_1 _21583_ (.A0(\digitop_pav2.ack_inst.buffer_ff[14] ),
    .A1(net1088),
    .S(net1160),
    .X(_01503_));
 mux2_1 _21584_ (.A0(\digitop_pav2.ack_inst.buffer_ff[15] ),
    .A1(net1085),
    .S(net1161),
    .X(_01504_));
 a41o_1 _21585_ (.A1(net1257),
    .A2(_08470_),
    .A3(_08474_),
    .A4(_09521_),
    .B1(\digitop_pav2.acc_activate ),
    .X(_01507_));
 and4_1 _21586_ (.A(_08050_),
    .B(_08060_),
    .C(_08062_),
    .D(_08084_),
    .X(_06147_));
 and3_1 _21587_ (.A(_08053_),
    .B(_08057_),
    .C(_06147_),
    .X(_06148_));
 or4_1 _21588_ (.A(_08058_),
    .B(_08073_),
    .C(_08077_),
    .D(_08080_),
    .X(_06149_));
 or4_1 _21589_ (.A(_08054_),
    .B(_08069_),
    .C(_08074_),
    .D(_08082_),
    .X(_06150_));
 and3_1 _21590_ (.A(_08064_),
    .B(_08067_),
    .C(_06148_),
    .X(_06151_));
 or3b_1 _21591_ (.A(_06149_),
    .B(_06150_),
    .C_N(_06151_),
    .X(_06152_));
 a41o_1 _21592_ (.A1(\digitop_pav2.access_inst.access_check0.ctrl_wcknzero_ck ),
    .A2(net1256),
    .A3(_07634_),
    .A4(_06152_),
    .B1(\digitop_pav2.access_inst.acc_wcknzero_o ),
    .X(_01516_));
 mux2_1 _21593_ (.A0(_08456_),
    .A1(\digitop_pav2.access_inst.access_check0.act_lock_st ),
    .S(_08038_),
    .X(_01518_));
 nand3_1 _21594_ (.A(\digitop_pav2.access_inst.access_ctrl0.crc_init_i ),
    .B(net1256),
    .C(\digitop_pav2.access_inst.access_ctrl0.crc_en_o ),
    .Y(_06153_));
 xor2_1 _21595_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[8] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[11] ),
    .X(_06154_));
 xnor2_2 _21596_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[0] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[4] ),
    .Y(_06155_));
 xnor2_1 _21597_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[12] ),
    .B(_06155_),
    .Y(_06156_));
 xnor2_1 _21598_ (.A(_06154_),
    .B(_06156_),
    .Y(_06157_));
 nand2_1 _21599_ (.A(net1019),
    .B(_06157_),
    .Y(_06158_));
 a221o_1 _21600_ (.A1(net811),
    .A2(_08044_),
    .B1(_08048_),
    .B2(net913),
    .C1(net964),
    .X(_06159_));
 nand2b_1 _21601_ (.A_N(_05267_),
    .B(net171),
    .Y(_06160_));
 xor2_1 _21602_ (.A(_06158_),
    .B(_06160_),
    .X(_06161_));
 a21oi_1 _21603_ (.A1(net1094),
    .A2(net962),
    .B1(_08045_),
    .Y(_06162_));
 a22o_2 _21604_ (.A1(net1035),
    .A2(net964),
    .B1(_08066_),
    .B2(_06162_),
    .X(_06163_));
 nand2_1 _21605_ (.A(net1107),
    .B(net170),
    .Y(_06164_));
 a21bo_1 _21606_ (.A1(net1097),
    .A2(net962),
    .B1_N(_08063_),
    .X(_06165_));
 o22ai_4 _21607_ (.A1(net1097),
    .A2(net963),
    .B1(_08045_),
    .B2(_06165_),
    .Y(_06166_));
 xnor2_2 _21608_ (.A(_06164_),
    .B(_06166_),
    .Y(_06167_));
 xor2_1 _21609_ (.A(_06163_),
    .B(_06167_),
    .X(_06168_));
 xnor2_1 _21610_ (.A(_06161_),
    .B(_06168_),
    .Y(_06169_));
 mux2_1 _21611_ (.A0(_06169_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[0] ),
    .S(net1029),
    .X(_01549_));
 nand2_1 _21612_ (.A(net1103),
    .B(net170),
    .Y(_06170_));
 nand2_1 _21613_ (.A(net1090),
    .B(net170),
    .Y(_06171_));
 mux2_1 _21614_ (.A0(net1090),
    .A1(_06171_),
    .S(_06170_),
    .X(_06172_));
 xnor2_2 _21615_ (.A(_06163_),
    .B(_06172_),
    .Y(_06173_));
 xor2_1 _21616_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[1] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[5] ),
    .X(_06174_));
 xor2_1 _21617_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[9] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[12] ),
    .X(_06175_));
 xnor2_1 _21618_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[13] ),
    .B(_06175_),
    .Y(_06176_));
 o21bai_1 _21619_ (.A1(_06174_),
    .A2(_06176_),
    .B1_N(\digitop_pav2.access_inst.access_ctrl0.crc_init_i ),
    .Y(_06177_));
 a21o_1 _21620_ (.A1(_06174_),
    .A2(_06176_),
    .B1(_06177_),
    .X(_06178_));
 nand2_1 _21621_ (.A(_05341_),
    .B(net170),
    .Y(_06179_));
 xnor2_1 _21622_ (.A(_06178_),
    .B(_06179_),
    .Y(_06180_));
 xnor2_1 _21623_ (.A(_06173_),
    .B(_06180_),
    .Y(_06181_));
 mux2_1 _21624_ (.A0(_06181_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[1] ),
    .S(net1028),
    .X(_01550_));
 nand2_1 _21625_ (.A(_05295_),
    .B(net170),
    .Y(_06182_));
 nand2_1 _21626_ (.A(_05296_),
    .B(net170),
    .Y(_06183_));
 xor2_1 _21627_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[10] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[13] ),
    .X(_06184_));
 xnor2_2 _21628_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[2] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[6] ),
    .Y(_06185_));
 xor2_1 _21629_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[14] ),
    .B(_06185_),
    .X(_06186_));
 a21oi_1 _21630_ (.A1(_06184_),
    .A2(_06186_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.crc_init_i ),
    .Y(_06187_));
 o21ai_1 _21631_ (.A1(_06184_),
    .A2(_06186_),
    .B1(_06187_),
    .Y(_06188_));
 xnor2_1 _21632_ (.A(_06183_),
    .B(_06188_),
    .Y(_06189_));
 mux2_1 _21633_ (.A0(_06189_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[2] ),
    .S(net1028),
    .X(_01551_));
 nand2_1 _21634_ (.A(_05301_),
    .B(net171),
    .Y(_06190_));
 xor2_1 _21635_ (.A(_06166_),
    .B(_06190_),
    .X(_06191_));
 xor2_2 _21636_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[3] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[7] ),
    .X(_06192_));
 xnor2_2 _21637_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[14] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[15] ),
    .Y(_06193_));
 xnor2_2 _21638_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[11] ),
    .B(_06193_),
    .Y(_06194_));
 xnor2_1 _21639_ (.A(_06192_),
    .B(_06194_),
    .Y(_06195_));
 nand2_1 _21640_ (.A(net1019),
    .B(_06195_),
    .Y(_06196_));
 xor2_1 _21641_ (.A(net1124),
    .B(net1113),
    .X(_06197_));
 nand2_1 _21642_ (.A(net171),
    .B(_06197_),
    .Y(_06198_));
 xor2_1 _21643_ (.A(_06196_),
    .B(_06198_),
    .X(_06199_));
 xnor2_1 _21644_ (.A(_06191_),
    .B(_06199_),
    .Y(_06200_));
 mux2_1 _21645_ (.A0(_06200_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[3] ),
    .S(net1029),
    .X(_01552_));
 and2b_1 _21646_ (.A_N(_05393_),
    .B(net171),
    .X(_06201_));
 xnor2_1 _21647_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[12] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[15] ),
    .Y(_06202_));
 xnor2_1 _21648_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[4] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[8] ),
    .Y(_06203_));
 o21ai_1 _21649_ (.A1(_06202_),
    .A2(_06203_),
    .B1(net1019),
    .Y(_06204_));
 a21o_1 _21650_ (.A1(_06202_),
    .A2(_06203_),
    .B1(_06204_),
    .X(_06205_));
 xnor2_1 _21651_ (.A(_06163_),
    .B(_06205_),
    .Y(_06206_));
 xnor2_1 _21652_ (.A(_06201_),
    .B(_06206_),
    .Y(_06207_));
 mux2_1 _21653_ (.A0(_06207_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[4] ),
    .S(net1029),
    .X(_01553_));
 xor2_1 _21654_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[5] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[8] ),
    .X(_06208_));
 xnor2_1 _21655_ (.A(_06155_),
    .B(_06208_),
    .Y(_06209_));
 xnor2_1 _21656_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[11] ),
    .B(_06176_),
    .Y(_06210_));
 o21ai_1 _21657_ (.A1(_06209_),
    .A2(_06210_),
    .B1(net1019),
    .Y(_06211_));
 a21o_1 _21658_ (.A1(_06209_),
    .A2(_06210_),
    .B1(_06211_),
    .X(_06212_));
 xnor2_1 _21659_ (.A(net1118),
    .B(_05267_),
    .Y(_06213_));
 nand2_1 _21660_ (.A(net171),
    .B(_06213_),
    .Y(_06214_));
 xnor2_1 _21661_ (.A(_06212_),
    .B(_06214_),
    .Y(_06215_));
 xnor2_1 _21662_ (.A(_06167_),
    .B(_06215_),
    .Y(_06216_));
 or2_1 _21663_ (.A(_06173_),
    .B(_06216_),
    .X(_06217_));
 a21oi_1 _21664_ (.A1(_06173_),
    .A2(_06216_),
    .B1(net1028),
    .Y(_06218_));
 a22o_1 _21665_ (.A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[5] ),
    .A2(net1028),
    .B1(_06217_),
    .B2(_06218_),
    .X(_01554_));
 nand2_1 _21666_ (.A(net1119),
    .B(net170),
    .Y(_06219_));
 nand2_1 _21667_ (.A(net1115),
    .B(net171),
    .Y(_06220_));
 a22o_1 _21668_ (.A1(net1118),
    .A2(net1115),
    .B1(_06219_),
    .B2(_06220_),
    .X(_06221_));
 nor2_1 _21669_ (.A(net1103),
    .B(_05294_),
    .Y(_06222_));
 and2_1 _21670_ (.A(net1103),
    .B(_05294_),
    .X(_06223_));
 o21a_1 _21671_ (.A1(_06222_),
    .A2(_06223_),
    .B1(net171),
    .X(_06224_));
 xor2_1 _21672_ (.A(_06221_),
    .B(_06224_),
    .X(_06225_));
 nand2_1 _21673_ (.A(net1131),
    .B(net170),
    .Y(_06226_));
 xnor2_1 _21674_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[13] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[14] ),
    .Y(_06227_));
 xnor2_1 _21675_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[12] ),
    .B(_06227_),
    .Y(_06228_));
 xnor2_1 _21676_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[6] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[10] ),
    .Y(_06229_));
 xnor2_1 _21677_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[9] ),
    .B(_06174_),
    .Y(_06230_));
 xnor2_1 _21678_ (.A(_06229_),
    .B(_06230_),
    .Y(_06231_));
 xnor2_1 _21679_ (.A(_06228_),
    .B(_06231_),
    .Y(_06232_));
 nand2_1 _21680_ (.A(net1019),
    .B(_06232_),
    .Y(_06233_));
 xor2_1 _21681_ (.A(_06163_),
    .B(_06233_),
    .X(_06234_));
 xnor2_1 _21682_ (.A(_06226_),
    .B(_06234_),
    .Y(_06235_));
 xnor2_1 _21683_ (.A(_06225_),
    .B(_06235_),
    .Y(_06236_));
 mux2_1 _21684_ (.A0(_06236_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[6] ),
    .S(net1028),
    .X(_01555_));
 nand2_2 _21685_ (.A(net1099),
    .B(net170),
    .Y(_06237_));
 xor2_2 _21686_ (.A(_06166_),
    .B(_06237_),
    .X(_06238_));
 xor2_1 _21687_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[7] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[10] ),
    .X(_06239_));
 xnor2_1 _21688_ (.A(_06185_),
    .B(_06239_),
    .Y(_06240_));
 xor2_1 _21689_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[13] ),
    .B(_06194_),
    .X(_06241_));
 o21ai_1 _21690_ (.A1(_06240_),
    .A2(_06241_),
    .B1(net1019),
    .Y(_06242_));
 a21o_1 _21691_ (.A1(_06240_),
    .A2(_06241_),
    .B1(_06242_),
    .X(_06243_));
 xnor2_1 _21692_ (.A(_06171_),
    .B(_06243_),
    .Y(_06244_));
 nand2_1 _21693_ (.A(net1128),
    .B(net1112),
    .Y(_06245_));
 or2_1 _21694_ (.A(net1128),
    .B(net1112),
    .X(_06246_));
 o22a_1 _21695_ (.A1(net1115),
    .A2(_06190_),
    .B1(_06220_),
    .B2(_05301_),
    .X(_06247_));
 xnor2_1 _21696_ (.A(_06244_),
    .B(_06247_),
    .Y(_06248_));
 and3_1 _21697_ (.A(net170),
    .B(_06245_),
    .C(_06246_),
    .X(_06249_));
 xor2_1 _21698_ (.A(_06238_),
    .B(_06249_),
    .X(_06250_));
 xnor2_1 _21699_ (.A(_06248_),
    .B(_06250_),
    .Y(_06251_));
 mux2_1 _21700_ (.A0(_06251_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[7] ),
    .S(net1028),
    .X(_01556_));
 xnor2_1 _21701_ (.A(_06190_),
    .B(_06198_),
    .Y(_06252_));
 xnor2_1 _21702_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[12] ),
    .B(_06193_),
    .Y(_06253_));
 xnor2_1 _21703_ (.A(_06154_),
    .B(_06192_),
    .Y(_06254_));
 a21oi_1 _21704_ (.A1(_06253_),
    .A2(_06254_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.crc_init_i ),
    .Y(_06255_));
 o21a_1 _21705_ (.A1(_06253_),
    .A2(_06254_),
    .B1(_06255_),
    .X(_06256_));
 xnor2_1 _21706_ (.A(_06252_),
    .B(_06256_),
    .Y(_06257_));
 xnor2_1 _21707_ (.A(_06168_),
    .B(_06257_),
    .Y(_06258_));
 mux2_1 _21708_ (.A0(_06258_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[8] ),
    .S(net1029),
    .X(_01557_));
 xor2_1 _21709_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[13] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[15] ),
    .X(_06259_));
 xnor2_1 _21710_ (.A(_06203_),
    .B(_06259_),
    .Y(_06260_));
 a21boi_1 _21711_ (.A1(_06175_),
    .A2(_06260_),
    .B1_N(net1019),
    .Y(_06261_));
 o21ai_1 _21712_ (.A1(_06175_),
    .A2(_06260_),
    .B1(_06261_),
    .Y(_06262_));
 xnor2_1 _21713_ (.A(_06201_),
    .B(_06262_),
    .Y(_06263_));
 xnor2_1 _21714_ (.A(_06173_),
    .B(_06263_),
    .Y(_06264_));
 mux2_1 _21715_ (.A0(_06264_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[9] ),
    .S(net1028),
    .X(_01558_));
 xor2_1 _21716_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[5] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[9] ),
    .X(_06265_));
 xnor2_1 _21717_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[14] ),
    .B(_06265_),
    .Y(_06266_));
 a21boi_1 _21718_ (.A1(_06184_),
    .A2(_06266_),
    .B1_N(net1019),
    .Y(_06267_));
 o21ai_1 _21719_ (.A1(_06184_),
    .A2(_06266_),
    .B1(_06267_),
    .Y(_06268_));
 xor2_1 _21720_ (.A(_06219_),
    .B(_06268_),
    .X(_06269_));
 xnor2_1 _21721_ (.A(_06224_),
    .B(_06269_),
    .Y(_06270_));
 mux2_1 _21722_ (.A0(_06270_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[10] ),
    .S(net1028),
    .X(_01559_));
 a21boi_1 _21723_ (.A1(_06194_),
    .A2(_06229_),
    .B1_N(_06153_),
    .Y(_06271_));
 o21ai_1 _21724_ (.A1(_06194_),
    .A2(_06229_),
    .B1(_06271_),
    .Y(_06272_));
 xor2_1 _21725_ (.A(_06237_),
    .B(_06272_),
    .X(_06273_));
 xnor2_1 _21726_ (.A(_06220_),
    .B(_06273_),
    .Y(_06274_));
 xnor2_1 _21727_ (.A(_06191_),
    .B(_06274_),
    .Y(_06275_));
 mux2_1 _21728_ (.A0(_06275_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[11] ),
    .S(net1029),
    .X(_01560_));
 nand2_1 _21729_ (.A(_05394_),
    .B(net171),
    .Y(_06276_));
 xnor2_1 _21730_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[8] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[15] ),
    .Y(_06277_));
 xnor2_1 _21731_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[7] ),
    .B(_06277_),
    .Y(_06278_));
 a21oi_1 _21732_ (.A1(_06155_),
    .A2(_06278_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.crc_init_i ),
    .Y(_06279_));
 o21ai_1 _21733_ (.A1(_06155_),
    .A2(_06278_),
    .B1(_06279_),
    .Y(_06280_));
 xnor2_1 _21734_ (.A(_06276_),
    .B(_06280_),
    .Y(_06281_));
 mux2_1 _21735_ (.A0(_06281_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[12] ),
    .S(net1029),
    .X(_01561_));
 a22o_1 _21736_ (.A1(net1107),
    .A2(net1103),
    .B1(_06164_),
    .B2(_06170_),
    .X(_06282_));
 xnor2_1 _21737_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[8] ),
    .B(_06230_),
    .Y(_06283_));
 nand2_1 _21738_ (.A(net1019),
    .B(_06283_),
    .Y(_06284_));
 xor2_1 _21739_ (.A(_06179_),
    .B(_06284_),
    .X(_06285_));
 xnor2_1 _21740_ (.A(_06282_),
    .B(_06285_),
    .Y(_06286_));
 mux2_1 _21741_ (.A0(_06286_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[13] ),
    .S(net1028),
    .X(_01562_));
 a22o_1 _21742_ (.A1(net1103),
    .A2(net1099),
    .B1(_06170_),
    .B2(_06237_),
    .X(_06287_));
 xor2_1 _21743_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[9] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[10] ),
    .X(_06288_));
 nand2_1 _21744_ (.A(_06185_),
    .B(_06288_),
    .Y(_06289_));
 or2_1 _21745_ (.A(_06185_),
    .B(_06288_),
    .X(_06290_));
 a21oi_1 _21746_ (.A1(_06289_),
    .A2(_06290_),
    .B1(\digitop_pav2.access_inst.access_ctrl0.crc_init_i ),
    .Y(_06291_));
 xnor2_1 _21747_ (.A(_06287_),
    .B(_06291_),
    .Y(_06292_));
 xnor2_1 _21748_ (.A(_06182_),
    .B(_06292_),
    .Y(_06293_));
 mux2_1 _21749_ (.A0(_06293_),
    .A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[14] ),
    .S(net1028),
    .X(_01563_));
 xor2_1 _21750_ (.A(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[10] ),
    .B(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[11] ),
    .X(_06294_));
 o21ai_1 _21751_ (.A1(_06192_),
    .A2(_06294_),
    .B1(net1019),
    .Y(_06295_));
 a21o_1 _21752_ (.A1(_06192_),
    .A2(_06294_),
    .B1(_06295_),
    .X(_06296_));
 xor2_1 _21753_ (.A(_06198_),
    .B(_06296_),
    .X(_06297_));
 nand2_1 _21754_ (.A(_06238_),
    .B(_06297_),
    .Y(_06298_));
 o21ba_1 _21755_ (.A1(_06238_),
    .A2(_06297_),
    .B1_N(net1029),
    .X(_06299_));
 a22o_1 _21756_ (.A1(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[15] ),
    .A2(net1029),
    .B1(_06298_),
    .B2(_06299_),
    .X(_01564_));
 and3_2 _21757_ (.A(_07031_),
    .B(net1143),
    .C(_07342_),
    .X(_06300_));
 nor2_1 _21758_ (.A(\digitop_pav2.access_inst.access_ctrl0.prev_busy ),
    .B(_02653_),
    .Y(_06301_));
 nor2_1 _21759_ (.A(_06300_),
    .B(_06301_),
    .Y(_06302_));
 nor2_1 _21760_ (.A(net1045),
    .B(_02653_),
    .Y(_06303_));
 nor2_1 _21761_ (.A(_06302_),
    .B(net677),
    .Y(_06304_));
 and3_1 _21762_ (.A(net1258),
    .B(_07524_),
    .C(net1016),
    .X(_06305_));
 nand2b_1 _21763_ (.A_N(_07525_),
    .B(net1016),
    .Y(_06306_));
 nand2_1 _21764_ (.A(_08324_),
    .B(net291),
    .Y(_06307_));
 and3_1 _21765_ (.A(_07383_),
    .B(_07393_),
    .C(_08909_),
    .X(_06308_));
 a31o_1 _21766_ (.A1(_07375_),
    .A2(_07405_),
    .A3(_08895_),
    .B1(_06308_),
    .X(_06309_));
 a211o_1 _21767_ (.A1(_07416_),
    .A2(_08908_),
    .B1(_06309_),
    .C1(_07394_),
    .X(_06310_));
 and3_1 _21768_ (.A(_07393_),
    .B(_07405_),
    .C(_08883_),
    .X(_06311_));
 a221o_1 _21769_ (.A1(_07385_),
    .A2(_08877_),
    .B1(_08889_),
    .B2(_07421_),
    .C1(_06311_),
    .X(_06312_));
 a2bb2o_1 _21770_ (.A1_N(_07402_),
    .A2_N(_08898_),
    .B1(_08900_),
    .B2(_07376_),
    .X(_06313_));
 a22o_1 _21771_ (.A1(_07422_),
    .A2(_08891_),
    .B1(_08911_),
    .B2(_07406_),
    .X(_06314_));
 and3_1 _21772_ (.A(_07375_),
    .B(_07383_),
    .C(_08890_),
    .X(_06315_));
 and3_1 _21773_ (.A(_07374_),
    .B(_07393_),
    .C(_08881_),
    .X(_06316_));
 a21o_1 _21774_ (.A1(_07415_),
    .A2(_08886_),
    .B1(_06316_),
    .X(_06317_));
 a211o_1 _21775_ (.A1(_07423_),
    .A2(_08913_),
    .B1(_06315_),
    .C1(_06317_),
    .X(_06318_));
 or4_1 _21776_ (.A(_06312_),
    .B(_06313_),
    .C(_06314_),
    .D(_06318_),
    .X(_06319_));
 a211o_1 _21777_ (.A1(_07420_),
    .A2(_08903_),
    .B1(_06310_),
    .C1(_06319_),
    .X(_06320_));
 nand2_1 _21778_ (.A(_07394_),
    .B(_08879_),
    .Y(_06321_));
 and3_1 _21779_ (.A(net1698),
    .B(_06320_),
    .C(_06321_),
    .X(_06322_));
 xor2_1 _21780_ (.A(net817),
    .B(_06322_),
    .X(_06323_));
 mux2_1 _21781_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[0] ),
    .A1(_06323_),
    .S(net807),
    .X(_06324_));
 nor2_1 _21782_ (.A(_06301_),
    .B(net676),
    .Y(_06325_));
 and2b_1 _21783_ (.A_N(net677),
    .B(_06302_),
    .X(_06326_));
 o211a_1 _21784_ (.A1(net291),
    .A2(_06324_),
    .B1(net570),
    .C1(_06307_),
    .X(_06327_));
 a31o_1 _21785_ (.A1(net1135),
    .A2(net181),
    .A3(_06304_),
    .B1(_06327_),
    .X(_06328_));
 a22o_1 _21786_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[0] ),
    .A2(net1201),
    .B1(net1010),
    .B2(_06328_),
    .X(_01568_));
 mux2_1 _21787_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[1] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[0] ),
    .S(net806),
    .X(_06329_));
 or2_1 _21788_ (.A(net290),
    .B(_06329_),
    .X(_06330_));
 o211a_1 _21789_ (.A1(_08293_),
    .A2(net254),
    .B1(net570),
    .C1(_06330_),
    .X(_06331_));
 a221o_1 _21790_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[0] ),
    .A2(net676),
    .B1(net571),
    .B2(_08056_),
    .C1(_06331_),
    .X(_06332_));
 a22o_1 _21791_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[1] ),
    .A2(net1200),
    .B1(net1009),
    .B2(_06332_),
    .X(_01569_));
 mux2_1 _21792_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[2] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[1] ),
    .S(net806),
    .X(_06333_));
 or2_1 _21793_ (.A(net290),
    .B(_06333_),
    .X(_06334_));
 o211a_1 _21794_ (.A1(_08259_),
    .A2(net254),
    .B1(net570),
    .C1(_06334_),
    .X(_06335_));
 a221o_1 _21795_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[1] ),
    .A2(net676),
    .B1(net571),
    .B2(_08058_),
    .C1(_06335_),
    .X(_06336_));
 a22o_1 _21796_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[2] ),
    .A2(net1203),
    .B1(net1009),
    .B2(_06336_),
    .X(_01570_));
 mux2_1 _21797_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[3] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[2] ),
    .S(net806),
    .X(_06337_));
 or2_1 _21798_ (.A(net290),
    .B(_06337_),
    .X(_06338_));
 o211a_1 _21799_ (.A1(_08153_),
    .A2(net254),
    .B1(net570),
    .C1(_06338_),
    .X(_06339_));
 a221o_1 _21800_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[2] ),
    .A2(net676),
    .B1(net571),
    .B2(_08077_),
    .C1(_06339_),
    .X(_06340_));
 a22o_1 _21801_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[3] ),
    .A2(net1200),
    .B1(net1009),
    .B2(_06340_),
    .X(_01571_));
 mux2_1 _21802_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[4] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[3] ),
    .S(net806),
    .X(_06341_));
 or2_1 _21803_ (.A(net290),
    .B(_06341_),
    .X(_06342_));
 o211a_1 _21804_ (.A1(_08171_),
    .A2(net254),
    .B1(net570),
    .C1(_06342_),
    .X(_06343_));
 a221o_1 _21805_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[3] ),
    .A2(net676),
    .B1(net571),
    .B2(_08080_),
    .C1(_06343_),
    .X(_06344_));
 a22o_1 _21806_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[4] ),
    .A2(net1203),
    .B1(net1009),
    .B2(_06344_),
    .X(_01572_));
 mux2_1 _21807_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[5] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[4] ),
    .S(net806),
    .X(_06345_));
 or2_1 _21808_ (.A(net290),
    .B(_06345_),
    .X(_06346_));
 o211a_1 _21809_ (.A1(_08372_),
    .A2(net254),
    .B1(net570),
    .C1(_06346_),
    .X(_06347_));
 a221o_1 _21810_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[4] ),
    .A2(net676),
    .B1(net571),
    .B2(_08052_),
    .C1(_06347_),
    .X(_06348_));
 a22o_1 _21811_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[5] ),
    .A2(net1200),
    .B1(net1009),
    .B2(_06348_),
    .X(_01573_));
 mux2_1 _21812_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[6] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[5] ),
    .S(net806),
    .X(_06349_));
 or2_1 _21813_ (.A(net290),
    .B(_06349_),
    .X(_06350_));
 o211a_1 _21814_ (.A1(_08225_),
    .A2(net254),
    .B1(net570),
    .C1(_06350_),
    .X(_06351_));
 a221o_1 _21815_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[5] ),
    .A2(net676),
    .B1(net571),
    .B2(_08082_),
    .C1(_06351_),
    .X(_06352_));
 a22o_1 _21816_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[6] ),
    .A2(net1200),
    .B1(net1009),
    .B2(_06352_),
    .X(_01574_));
 nor2_1 _21817_ (.A(_08341_),
    .B(net254),
    .Y(_06353_));
 mux2_1 _21818_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[7] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[6] ),
    .S(net806),
    .X(_06354_));
 a211o_1 _21819_ (.A1(net254),
    .A2(_06354_),
    .B1(_06353_),
    .C1(_06300_),
    .X(_06355_));
 nand2_1 _21820_ (.A(_08055_),
    .B(_06300_),
    .Y(_06356_));
 a32o_1 _21821_ (.A1(net1044),
    .A2(_08054_),
    .A3(_06301_),
    .B1(net676),
    .B2(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[6] ),
    .X(_06357_));
 a31o_1 _21822_ (.A1(_06325_),
    .A2(_06355_),
    .A3(_06356_),
    .B1(_06357_),
    .X(_06358_));
 a22o_1 _21823_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[7] ),
    .A2(net1200),
    .B1(net1009),
    .B2(_06358_),
    .X(_01575_));
 mux2_1 _21824_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[8] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[7] ),
    .S(net806),
    .X(_06359_));
 mux2_1 _21825_ (.A0(_08356_),
    .A1(_06359_),
    .S(net254),
    .X(_06360_));
 mux2_1 _21826_ (.A0(_06360_),
    .A1(_08069_),
    .S(_06300_),
    .X(_06361_));
 a22o_1 _21827_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[7] ),
    .A2(net676),
    .B1(_06325_),
    .B2(_06361_),
    .X(_06362_));
 a31o_1 _21828_ (.A1(net1044),
    .A2(_08069_),
    .A3(_06301_),
    .B1(_06362_),
    .X(_06363_));
 a22o_1 _21829_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[8] ),
    .A2(net1200),
    .B1(net1009),
    .B2(_06363_),
    .X(_01576_));
 mux2_1 _21830_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[9] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[8] ),
    .S(net806),
    .X(_06364_));
 or2_1 _21831_ (.A(net290),
    .B(_06364_),
    .X(_06365_));
 o211a_1 _21832_ (.A1(_08188_),
    .A2(net254),
    .B1(net570),
    .C1(_06365_),
    .X(_06366_));
 a221o_1 _21833_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[8] ),
    .A2(net676),
    .B1(net571),
    .B2(_08061_),
    .C1(_06366_),
    .X(_06367_));
 a22o_1 _21834_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[9] ),
    .A2(net1200),
    .B1(net1009),
    .B2(_06367_),
    .X(_01577_));
 mux2_1 _21835_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[10] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[9] ),
    .S(net806),
    .X(_06368_));
 or2_1 _21836_ (.A(net290),
    .B(_06368_),
    .X(_06369_));
 o211a_1 _21837_ (.A1(_08276_),
    .A2(net255),
    .B1(net570),
    .C1(_06369_),
    .X(_06370_));
 a221o_1 _21838_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[9] ),
    .A2(net677),
    .B1(net571),
    .B2(_08074_),
    .C1(_06370_),
    .X(_06371_));
 a22o_1 _21839_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[10] ),
    .A2(net1200),
    .B1(net1009),
    .B2(_06371_),
    .X(_01578_));
 mux2_1 _21840_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[11] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[10] ),
    .S(net807),
    .X(_06372_));
 or2_1 _21841_ (.A(net290),
    .B(_06372_),
    .X(_06373_));
 o211a_1 _21842_ (.A1(_08387_),
    .A2(net255),
    .B1(_06326_),
    .C1(_06373_),
    .X(_06374_));
 a221o_1 _21843_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[10] ),
    .A2(net677),
    .B1(net571),
    .B2(_08065_),
    .C1(_06374_),
    .X(_06375_));
 a22o_1 _21844_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[11] ),
    .A2(net1200),
    .B1(net1010),
    .B2(_06375_),
    .X(_01579_));
 mux2_1 _21845_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[12] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[11] ),
    .S(net807),
    .X(_06376_));
 or2_1 _21846_ (.A(net291),
    .B(_06376_),
    .X(_06377_));
 o211a_1 _21847_ (.A1(_08308_),
    .A2(net255),
    .B1(_06326_),
    .C1(_06377_),
    .X(_06378_));
 a221o_1 _21848_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[11] ),
    .A2(net677),
    .B1(_06304_),
    .B2(_08068_),
    .C1(_06378_),
    .X(_06379_));
 a22o_1 _21849_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[12] ),
    .A2(net1200),
    .B1(net1010),
    .B2(_06379_),
    .X(_01580_));
 mux2_1 _21850_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[13] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[12] ),
    .S(net807),
    .X(_06380_));
 or2_1 _21851_ (.A(net290),
    .B(_06380_),
    .X(_06381_));
 o211a_1 _21852_ (.A1(_08207_),
    .A2(net255),
    .B1(_06326_),
    .C1(_06381_),
    .X(_06382_));
 a221o_1 _21853_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[12] ),
    .A2(net677),
    .B1(net571),
    .B2(_08073_),
    .C1(_06382_),
    .X(_06383_));
 a22o_1 _21854_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[13] ),
    .A2(net1203),
    .B1(net1010),
    .B2(_06383_),
    .X(_01581_));
 mux2_1 _21855_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[14] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[13] ),
    .S(net807),
    .X(_06384_));
 or2_1 _21856_ (.A(net291),
    .B(_06384_),
    .X(_06385_));
 o211a_1 _21857_ (.A1(_08399_),
    .A2(net255),
    .B1(_06326_),
    .C1(_06385_),
    .X(_06386_));
 a221o_1 _21858_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[13] ),
    .A2(net677),
    .B1(_06304_),
    .B2(_08085_),
    .C1(_06386_),
    .X(_06387_));
 a22o_1 _21859_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[14] ),
    .A2(net1202),
    .B1(net1010),
    .B2(_06387_),
    .X(_01582_));
 mux2_1 _21860_ (.A0(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[15] ),
    .A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[14] ),
    .S(net807),
    .X(_06388_));
 or2_1 _21861_ (.A(net291),
    .B(_06388_),
    .X(_06389_));
 o211a_1 _21862_ (.A1(_08241_),
    .A2(net255),
    .B1(net570),
    .C1(_06389_),
    .X(_06390_));
 a221o_1 _21863_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[14] ),
    .A2(net677),
    .B1(_06304_),
    .B2(_08051_),
    .C1(_06390_),
    .X(_06391_));
 a22o_1 _21864_ (.A1(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[15] ),
    .A2(net1202),
    .B1(net1010),
    .B2(_06391_),
    .X(_01583_));
 mux2_1 _21865_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt0_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[0] ),
    .S(net151),
    .X(_01585_));
 mux2_1 _21866_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt1_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[1] ),
    .S(net151),
    .X(_01586_));
 mux2_1 _21867_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt2_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[2] ),
    .S(net151),
    .X(_01587_));
 mux2_1 _21868_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt3_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[3] ),
    .S(net151),
    .X(_01588_));
 mux2_1 _21869_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt4_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[4] ),
    .S(net151),
    .X(_01589_));
 mux2_1 _21870_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt5_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[5] ),
    .S(net151),
    .X(_01590_));
 mux2_1 _21871_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt6_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[6] ),
    .S(net152),
    .X(_01591_));
 mux2_1 _21872_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt7_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[7] ),
    .S(net152),
    .X(_01592_));
 mux2_1 _21873_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt8_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[8] ),
    .S(net152),
    .X(_01593_));
 mux2_1 _21874_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt9_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[9] ),
    .S(net151),
    .X(_01594_));
 mux2_1 _21875_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt10_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[10] ),
    .S(net152),
    .X(_01595_));
 mux2_1 _21876_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt11_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[11] ),
    .S(net151),
    .X(_01596_));
 mux2_1 _21877_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt12_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[12] ),
    .S(net152),
    .X(_01597_));
 mux2_1 _21878_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt13_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[13] ),
    .S(net151),
    .X(_01598_));
 mux2_1 _21879_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt14_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[14] ),
    .S(net152),
    .X(_01599_));
 mux2_1 _21880_ (.A0(\digitop_pav2.stadly_memctrl_wr_dt15_1.Y ),
    .A1(\digitop_pav2.memctrl_inst.flops_0x081[15] ),
    .S(net152),
    .X(_01600_));
 nor2_1 _21881_ (.A(_10992_),
    .B(_11003_),
    .Y(_06392_));
 o22a_1 _21882_ (.A1(\digitop_pav2.pie_inst.fsm.state[0] ),
    .A2(_10981_),
    .B1(_10990_),
    .B2(_06392_),
    .X(_06393_));
 or2_1 _21883_ (.A(\digitop_pav2.pie_inst.fsm.pivot[5] ),
    .B(net495),
    .X(_06394_));
 a211o_1 _21884_ (.A1(\digitop_pav2.pie_inst.fsm.past_ctr[1] ),
    .A2(\digitop_pav2.pie_inst.fsm.pivot[1] ),
    .B1(\digitop_pav2.pie_inst.fsm.pivot[0] ),
    .C1(_07146_),
    .X(_06395_));
 o221a_1 _21885_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[2] ),
    .A2(_09576_),
    .B1(_10957_),
    .B2(\digitop_pav2.pie_inst.fsm.pivot[1] ),
    .C1(_06395_),
    .X(_06396_));
 a221o_1 _21886_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[2] ),
    .A2(_09576_),
    .B1(_09583_),
    .B2(net1301),
    .C1(_06396_),
    .X(_06397_));
 o221a_1 _21887_ (.A1(net1301),
    .A2(_09583_),
    .B1(_10949_),
    .B2(\digitop_pav2.pie_inst.fsm.pivot[4] ),
    .C1(_06397_),
    .X(_06398_));
 a221o_1 _21888_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[5] ),
    .A2(net495),
    .B1(_10949_),
    .B2(\digitop_pav2.pie_inst.fsm.pivot[4] ),
    .C1(_06398_),
    .X(_06399_));
 a22o_1 _21889_ (.A1(net1300),
    .A2(net493),
    .B1(_06394_),
    .B2(_06399_),
    .X(_06400_));
 o221a_1 _21890_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[7] ),
    .A2(net494),
    .B1(net493),
    .B2(net1300),
    .C1(_06400_),
    .X(_06401_));
 a221o_1 _21891_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[7] ),
    .A2(net494),
    .B1(net491),
    .B2(\digitop_pav2.pie_inst.fsm.pivot[8] ),
    .C1(_06401_),
    .X(_06402_));
 o21ai_1 _21892_ (.A1(\digitop_pav2.pie_inst.fsm.pivot[8] ),
    .A2(net491),
    .B1(_06402_),
    .Y(_06403_));
 o211a_1 _21893_ (.A1(\digitop_pav2.pie_inst.fsm.dif_pos_fix[9] ),
    .A2(_06403_),
    .B1(_11004_),
    .C1(_10981_),
    .X(_06404_));
 mux2_1 _21894_ (.A0(_06404_),
    .A1(\digitop_pav2.crc_inst.dt_rx_i ),
    .S(_06393_),
    .X(_01601_));
 or2_1 _21895_ (.A(net1456),
    .B(\digitop_pav2.sync_inst.inst_rstx.gray_counter[1] ),
    .X(_06405_));
 mux2_1 _21896_ (.A0(_07236_),
    .A1(\digitop_pav2.sync_inst.inst_rstx.gray_counter[0] ),
    .S(_06405_),
    .X(_01606_));
 mux2_1 _21897_ (.A0(\digitop_pav2.proc_ctrl_inst.ebv.state[14] ),
    .A1(\digitop_pav2.proc_ctrl_inst.ebv.state[12] ),
    .S(net971),
    .X(_01607_));
 mux2_1 _21898_ (.A0(\digitop_pav2.proc_ctrl_inst.ebv.state[13] ),
    .A1(\digitop_pav2.proc_ctrl_inst.ebv.state[11] ),
    .S(net970),
    .X(_01608_));
 mux2_1 _21899_ (.A0(\digitop_pav2.proc_ctrl_inst.ebv.state[12] ),
    .A1(\digitop_pav2.proc_ctrl_inst.ebv.state[5] ),
    .S(net970),
    .X(_01609_));
 mux2_1 _21900_ (.A0(\digitop_pav2.proc_ctrl_inst.ebv.state[11] ),
    .A1(\digitop_pav2.proc_ctrl_inst.ebv.state[8] ),
    .S(net970),
    .X(_01610_));
 mux2_1 _21901_ (.A0(\digitop_pav2.proc_ctrl_inst.ebv.state[10] ),
    .A1(\digitop_pav2.proc_ctrl_inst.ebv.state[14] ),
    .S(net971),
    .X(_01611_));
 mux2_1 _21902_ (.A0(\digitop_pav2.proc_ctrl_inst.ebv.state[9] ),
    .A1(\digitop_pav2.proc_ctrl_inst.ebv.state[10] ),
    .S(net971),
    .X(_01612_));
 mux2_1 _21903_ (.A0(\digitop_pav2.proc_ctrl_inst.ebv.state[7] ),
    .A1(\digitop_pav2.proc_ctrl_inst.ebv.state[6] ),
    .S(net970),
    .X(_01613_));
 mux2_1 _21904_ (.A0(\digitop_pav2.proc_ctrl_inst.ebv.state[6] ),
    .A1(\digitop_pav2.proc_ctrl_inst.ebv.state[13] ),
    .S(net970),
    .X(_01614_));
 mux2_1 _21905_ (.A0(\digitop_pav2.proc_ctrl_inst.ebv.state[5] ),
    .A1(\digitop_pav2.proc_ctrl_inst.ebv.state[4] ),
    .S(net970),
    .X(_01615_));
 mux2_1 _21906_ (.A0(\digitop_pav2.proc_ctrl_inst.ebv.state[3] ),
    .A1(\digitop_pav2.proc_ctrl_inst.ebv.state[7] ),
    .S(net971),
    .X(_01616_));
 mux2_1 _21907_ (.A0(\digitop_pav2.proc_ctrl_inst.ebv.state[2] ),
    .A1(\digitop_pav2.proc_ctrl_inst.ebv.state[9] ),
    .S(net971),
    .X(_01617_));
 mux2_1 _21908_ (.A0(\digitop_pav2.proc_ctrl_inst.ebv.state[1] ),
    .A1(\digitop_pav2.proc_ctrl_inst.ebv.state[3] ),
    .S(net971),
    .X(_01618_));
 o21a_1 _21909_ (.A1(\digitop_pav2.proc_ctrl_inst.ebv.state[2] ),
    .A2(\digitop_pav2.proc_ctrl_inst.ebv.state[1] ),
    .B1(net970),
    .X(_06406_));
 a21o_1 _21910_ (.A1(_07111_),
    .A2(\digitop_pav2.proc_ctrl_inst.ebv.state[0] ),
    .B1(_06406_),
    .X(_01619_));
 mux2_1 _21911_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[15] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[11] ),
    .S(net1167),
    .X(_01620_));
 mux2_1 _21912_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[14] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[6] ),
    .S(net1166),
    .X(_01621_));
 mux2_1 _21913_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[13] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[5] ),
    .S(net1166),
    .X(_01622_));
 mux2_1 _21914_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[12] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[8] ),
    .S(net1167),
    .X(_01623_));
 mux2_1 _21915_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[11] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[3] ),
    .S(net1166),
    .X(_01624_));
 mux2_1 _21916_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[10] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[14] ),
    .S(net1166),
    .X(_01625_));
 mux2_1 _21917_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[9] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[13] ),
    .S(net1167),
    .X(_01626_));
 mux2_1 _21918_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[8] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[0] ),
    .S(net1167),
    .X(_01627_));
 mux2_1 _21919_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[7] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[15] ),
    .S(net1166),
    .X(_01628_));
 mux2_1 _21920_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[6] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[4] ),
    .S(net1166),
    .X(_01629_));
 mux2_1 _21921_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[5] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[7] ),
    .S(net1166),
    .X(_01630_));
 mux2_1 _21922_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[4] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[12] ),
    .S(net1166),
    .X(_01631_));
 mux2_1 _21923_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[3] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[2] ),
    .S(net1166),
    .X(_01632_));
 mux2_1 _21924_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[2] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[10] ),
    .S(net1166),
    .X(_01633_));
 mux2_1 _21925_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[1] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[9] ),
    .S(net1167),
    .X(_01634_));
 mux2_1 _21926_ (.A0(\digitop_pav2.proc_ctrl_inst.inst_checker.state[0] ),
    .A1(\digitop_pav2.proc_ctrl_inst.inst_checker.state[1] ),
    .S(net1167),
    .X(_01635_));
 mux2_1 _21927_ (.A0(\digitop_pav2.sec_inst.ld_mem.st[3] ),
    .A1(\digitop_pav2.sec_inst.ld_mem.st[0] ),
    .S(_09660_),
    .X(_01636_));
 mux2_1 _21928_ (.A0(\digitop_pav2.sec_inst.ld_mem.st[2] ),
    .A1(\digitop_pav2.sec_inst.ld_mem.st[3] ),
    .S(_09660_),
    .X(_01637_));
 mux2_1 _21929_ (.A0(net707),
    .A1(net701),
    .S(_08504_),
    .X(_01638_));
 mux2_1 _21930_ (.A0(_04377_),
    .A1(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[1] ),
    .S(_09615_),
    .X(_01639_));
 nor2_2 _21931_ (.A(net84),
    .B(net86),
    .Y(_06407_));
 or2_2 _21932_ (.A(net84),
    .B(net86),
    .X(_06408_));
 nand2_1 _21933_ (.A(net94),
    .B(net953),
    .Y(_06409_));
 or2_2 _21934_ (.A(net907),
    .B(_06409_),
    .X(_06410_));
 o21ai_4 _21935_ (.A1(\stadly_mpw03_prog_rise_9.Y ),
    .A2(net1327),
    .B1(_09416_),
    .Y(_06411_));
 or4_1 _21936_ (.A(net778),
    .B(net618),
    .C(_06410_),
    .D(net867),
    .X(_06412_));
 mux2_1 _21937_ (.A0(net1358),
    .A1(\vmem[511] ),
    .S(_06412_),
    .X(_01640_));
 nand2_1 _21938_ (.A(net93),
    .B(net953),
    .Y(_06413_));
 or2_2 _21939_ (.A(net907),
    .B(_06413_),
    .X(_06414_));
 or4_1 _21940_ (.A(net783),
    .B(net623),
    .C(net871),
    .D(_06414_),
    .X(_06415_));
 mux2_1 _21941_ (.A0(net1368),
    .A1(\vmem[510] ),
    .S(_06415_),
    .X(_01641_));
 nor2_1 _21942_ (.A(_10836_),
    .B(net934),
    .Y(_06416_));
 nand2_2 _21943_ (.A(net897),
    .B(_06416_),
    .Y(_06417_));
 or4_1 _21944_ (.A(net774),
    .B(net616),
    .C(net865),
    .D(_06417_),
    .X(_06418_));
 mux2_1 _21945_ (.A0(net1353),
    .A1(\vmem[509] ),
    .S(_06418_),
    .X(_01642_));
 nand2_1 _21946_ (.A(net91),
    .B(net953),
    .Y(_06419_));
 or2_2 _21947_ (.A(net909),
    .B(_06419_),
    .X(_06420_));
 or4_1 _21948_ (.A(net796),
    .B(net635),
    .C(net881),
    .D(_06420_),
    .X(_06421_));
 mux2_1 _21949_ (.A0(net1387),
    .A1(\vmem[508] ),
    .S(_06421_),
    .X(_01643_));
 nor2_1 _21950_ (.A(_10835_),
    .B(net932),
    .Y(_06422_));
 nand2_2 _21951_ (.A(net899),
    .B(_06422_),
    .Y(_06423_));
 or4_1 _21952_ (.A(net779),
    .B(net620),
    .C(net868),
    .D(_06423_),
    .X(_06424_));
 mux2_1 _21953_ (.A0(net1361),
    .A1(\vmem[507] ),
    .S(_06424_),
    .X(_01644_));
 nand2_1 _21954_ (.A(net89),
    .B(net953),
    .Y(_06425_));
 or2_2 _21955_ (.A(net908),
    .B(_06425_),
    .X(_06426_));
 or4_1 _21956_ (.A(net771),
    .B(net614),
    .C(net858),
    .D(_06426_),
    .X(_06427_));
 mux2_1 _21957_ (.A0(net1346),
    .A1(\vmem[506] ),
    .S(_06427_),
    .X(_01645_));
 nor2_1 _21958_ (.A(_10834_),
    .B(net939),
    .Y(_06428_));
 nand2_2 _21959_ (.A(net900),
    .B(_06428_),
    .Y(_06429_));
 or4_1 _21960_ (.A(net788),
    .B(net625),
    .C(net874),
    .D(_06429_),
    .X(_06430_));
 mux2_1 _21961_ (.A0(net1372),
    .A1(\vmem[505] ),
    .S(_06430_),
    .X(_01646_));
 nor2_1 _21962_ (.A(_10833_),
    .B(net920),
    .Y(_06431_));
 nand2_2 _21963_ (.A(net890),
    .B(_06431_),
    .Y(_06432_));
 or4_1 _21964_ (.A(net764),
    .B(net610),
    .C(net857),
    .D(_06432_),
    .X(_06433_));
 mux2_1 _21965_ (.A0(net1337),
    .A1(\vmem[504] ),
    .S(_06433_),
    .X(_01647_));
 nand2_1 _21966_ (.A(net101),
    .B(net953),
    .Y(_06434_));
 or2_2 _21967_ (.A(net908),
    .B(_06434_),
    .X(_06435_));
 or4_1 _21968_ (.A(net774),
    .B(net616),
    .C(net864),
    .D(_06435_),
    .X(_06436_));
 mux2_1 _21969_ (.A0(net1352),
    .A1(\vmem[503] ),
    .S(_06436_),
    .X(_01648_));
 nand2_1 _21970_ (.A(net100),
    .B(net953),
    .Y(_06437_));
 or2_2 _21971_ (.A(net909),
    .B(_06437_),
    .X(_06438_));
 or4_1 _21972_ (.A(net797),
    .B(net637),
    .C(net883),
    .D(_06438_),
    .X(_06439_));
 mux2_1 _21973_ (.A0(net1390),
    .A1(\vmem[502] ),
    .S(_06439_),
    .X(_01649_));
 nor2_1 _21974_ (.A(_10830_),
    .B(net917),
    .Y(_06440_));
 nand2_2 _21975_ (.A(net887),
    .B(_06440_),
    .Y(_06441_));
 or4_1 _21976_ (.A(net762),
    .B(net607),
    .C(net856),
    .D(_06441_),
    .X(_06442_));
 mux2_1 _21977_ (.A0(net1334),
    .A1(\vmem[501] ),
    .S(_06442_),
    .X(_01650_));
 nand2_1 _21978_ (.A(net98),
    .B(net954),
    .Y(_06443_));
 or2_2 _21979_ (.A(net909),
    .B(_06443_),
    .X(_06444_));
 or4_1 _21980_ (.A(net792),
    .B(net630),
    .C(net880),
    .D(_06444_),
    .X(_06445_));
 mux2_1 _21981_ (.A0(net1380),
    .A1(\vmem[500] ),
    .S(_06445_),
    .X(_01651_));
 nor2_1 _21982_ (.A(_10829_),
    .B(net917),
    .Y(_06446_));
 nand2_2 _21983_ (.A(net888),
    .B(_06446_),
    .Y(_06447_));
 or4_1 _21984_ (.A(net758),
    .B(net604),
    .C(net853),
    .D(_06447_),
    .X(_06448_));
 mux2_1 _21985_ (.A0(net1328),
    .A1(\vmem[499] ),
    .S(_06448_),
    .X(_01652_));
 nand2_1 _21986_ (.A(net96),
    .B(net954),
    .Y(_06449_));
 or2_2 _21987_ (.A(net909),
    .B(_06449_),
    .X(_06450_));
 or4_1 _21988_ (.A(net792),
    .B(net633),
    .C(net880),
    .D(_06450_),
    .X(_06451_));
 mux2_1 _21989_ (.A0(net1381),
    .A1(\vmem[498] ),
    .S(_06451_),
    .X(_01653_));
 nor2_1 _21990_ (.A(_10826_),
    .B(net940),
    .Y(_06452_));
 nand2_2 _21991_ (.A(net900),
    .B(_06452_),
    .Y(_06453_));
 or4_1 _21992_ (.A(net789),
    .B(net628),
    .C(net878),
    .D(_06453_),
    .X(_06454_));
 mux2_1 _21993_ (.A0(net1377),
    .A1(\vmem[497] ),
    .S(_06454_),
    .X(_01654_));
 o21a_1 _21994_ (.A1(_10819_),
    .A2(_10822_),
    .B1(_10821_),
    .X(_06455_));
 nor2_1 _21995_ (.A(net923),
    .B(_06455_),
    .Y(_06456_));
 nand2_2 _21996_ (.A(net892),
    .B(_06456_),
    .Y(_06457_));
 or4_1 _21997_ (.A(net767),
    .B(net613),
    .C(net859),
    .D(_06457_),
    .X(_06458_));
 mux2_1 _21998_ (.A0(net1342),
    .A1(\vmem[496] ),
    .S(_06458_),
    .X(_01655_));
 nand2_1 _21999_ (.A(net94),
    .B(net931),
    .Y(_06459_));
 or2_2 _22000_ (.A(net907),
    .B(_06459_),
    .X(_06460_));
 or4_1 _22001_ (.A(net777),
    .B(net619),
    .C(net866),
    .D(_06460_),
    .X(_06461_));
 mux2_1 _22002_ (.A0(net1356),
    .A1(\vmem[495] ),
    .S(_06461_),
    .X(_01656_));
 nand2_1 _22003_ (.A(net93),
    .B(net935),
    .Y(_06462_));
 or2_2 _22004_ (.A(net907),
    .B(_06462_),
    .X(_06463_));
 or4_1 _22005_ (.A(net793),
    .B(net632),
    .C(net879),
    .D(_06463_),
    .X(_06464_));
 mux2_1 _22006_ (.A0(net1369),
    .A1(\vmem[494] ),
    .S(_06464_),
    .X(_01657_));
 nor2_1 _22007_ (.A(_10836_),
    .B(net953),
    .Y(_06465_));
 nand2_2 _22008_ (.A(net897),
    .B(_06465_),
    .Y(_06466_));
 or4_1 _22009_ (.A(net784),
    .B(net621),
    .C(net872),
    .D(_06466_),
    .X(_06467_));
 mux2_1 _22010_ (.A0(net1365),
    .A1(\vmem[493] ),
    .S(_06467_),
    .X(_01658_));
 nand2_1 _22011_ (.A(net91),
    .B(net942),
    .Y(_06468_));
 or2_2 _22012_ (.A(net909),
    .B(_06468_),
    .X(_06469_));
 or4_1 _22013_ (.A(net796),
    .B(net634),
    .C(net877),
    .D(_06469_),
    .X(_06470_));
 mux2_1 _22014_ (.A0(net1386),
    .A1(\vmem[492] ),
    .S(_06470_),
    .X(_01659_));
 nor2_1 _22015_ (.A(_10835_),
    .B(net953),
    .Y(_06471_));
 nand2_2 _22016_ (.A(net896),
    .B(_06471_),
    .Y(_06472_));
 or4_1 _22017_ (.A(net779),
    .B(net620),
    .C(net868),
    .D(_06472_),
    .X(_06473_));
 mux2_1 _22018_ (.A0(net1361),
    .A1(\vmem[491] ),
    .S(_06473_),
    .X(_01660_));
 nand2_1 _22019_ (.A(net89),
    .B(net927),
    .Y(_06474_));
 or2_2 _22020_ (.A(net908),
    .B(_06474_),
    .X(_06475_));
 or4_1 _22021_ (.A(net771),
    .B(net614),
    .C(net858),
    .D(_06475_),
    .X(_06476_));
 mux2_1 _22022_ (.A0(net1346),
    .A1(\vmem[490] ),
    .S(_06476_),
    .X(_01661_));
 nor2_1 _22023_ (.A(_10834_),
    .B(net954),
    .Y(_06477_));
 nand2_2 _22024_ (.A(net900),
    .B(_06477_),
    .Y(_06478_));
 or4_1 _22025_ (.A(net788),
    .B(net626),
    .C(net876),
    .D(_06478_),
    .X(_06479_));
 mux2_1 _22026_ (.A0(net1374),
    .A1(\vmem[489] ),
    .S(_06479_),
    .X(_01662_));
 nor2_1 _22027_ (.A(_10833_),
    .B(net952),
    .Y(_06480_));
 nand2_2 _22028_ (.A(net890),
    .B(_06480_),
    .Y(_06481_));
 or4_1 _22029_ (.A(net764),
    .B(net610),
    .C(net854),
    .D(_06481_),
    .X(_06482_));
 mux2_1 _22030_ (.A0(net1336),
    .A1(\vmem[488] ),
    .S(_06482_),
    .X(_01663_));
 nand2_1 _22031_ (.A(net101),
    .B(net928),
    .Y(_06483_));
 or2_2 _22032_ (.A(net908),
    .B(_06483_),
    .X(_06484_));
 or4_1 _22033_ (.A(net774),
    .B(net616),
    .C(net864),
    .D(_06484_),
    .X(_06485_));
 mux2_1 _22034_ (.A0(net1354),
    .A1(\vmem[487] ),
    .S(_06485_),
    .X(_01664_));
 nand2_1 _22035_ (.A(net100),
    .B(net948),
    .Y(_06486_));
 or2_2 _22036_ (.A(net909),
    .B(_06486_),
    .X(_06487_));
 or4_1 _22037_ (.A(net797),
    .B(net636),
    .C(net883),
    .D(_06487_),
    .X(_06488_));
 mux2_1 _22038_ (.A0(net1390),
    .A1(\vmem[486] ),
    .S(_06488_),
    .X(_01665_));
 nor2_1 _22039_ (.A(_10830_),
    .B(net952),
    .Y(_06489_));
 nand2_2 _22040_ (.A(net889),
    .B(_06489_),
    .Y(_06490_));
 or4_1 _22041_ (.A(net762),
    .B(net607),
    .C(_06411_),
    .D(_06490_),
    .X(_06491_));
 mux2_1 _22042_ (.A0(net1334),
    .A1(\vmem[485] ),
    .S(_06491_),
    .X(_01666_));
 nand2_1 _22043_ (.A(net98),
    .B(net944),
    .Y(_06492_));
 or2_2 _22044_ (.A(net909),
    .B(_06492_),
    .X(_06493_));
 or4_1 _22045_ (.A(net792),
    .B(net630),
    .C(net880),
    .D(_06493_),
    .X(_06494_));
 mux2_1 _22046_ (.A0(net1380),
    .A1(\vmem[484] ),
    .S(_06494_),
    .X(_01667_));
 nor2_1 _22047_ (.A(_10829_),
    .B(net952),
    .Y(_06495_));
 nand2_2 _22048_ (.A(net887),
    .B(_06495_),
    .Y(_06496_));
 or4_1 _22049_ (.A(net758),
    .B(net604),
    .C(net853),
    .D(_06496_),
    .X(_06497_));
 mux2_1 _22050_ (.A0(net1328),
    .A1(\vmem[483] ),
    .S(_06497_),
    .X(_01668_));
 nand2_1 _22051_ (.A(net96),
    .B(net940),
    .Y(_06498_));
 or2_2 _22052_ (.A(net909),
    .B(_06498_),
    .X(_06499_));
 or4_1 _22053_ (.A(net795),
    .B(net633),
    .C(net876),
    .D(_06499_),
    .X(_06500_));
 mux2_1 _22054_ (.A0(net1381),
    .A1(\vmem[482] ),
    .S(_06500_),
    .X(_01669_));
 nor2_1 _22055_ (.A(_10826_),
    .B(net954),
    .Y(_06501_));
 nand2_2 _22056_ (.A(net901),
    .B(_06501_),
    .Y(_06502_));
 or4_1 _22057_ (.A(net789),
    .B(net627),
    .C(net877),
    .D(_06502_),
    .X(_06503_));
 mux2_1 _22058_ (.A0(net1377),
    .A1(\vmem[481] ),
    .S(_06503_),
    .X(_01670_));
 nor2_1 _22059_ (.A(net952),
    .B(_06455_),
    .Y(_06504_));
 nand2_2 _22060_ (.A(net892),
    .B(_06504_),
    .Y(_06505_));
 or4_1 _22061_ (.A(net766),
    .B(net613),
    .C(net860),
    .D(_06505_),
    .X(_06506_));
 mux2_1 _22062_ (.A0(net1342),
    .A1(\vmem[480] ),
    .S(_06506_),
    .X(_01671_));
 or2_2 _22063_ (.A(net896),
    .B(_06409_),
    .X(_06507_));
 or4_1 _22064_ (.A(net777),
    .B(net618),
    .C(net867),
    .D(_06507_),
    .X(_06508_));
 mux2_1 _22065_ (.A0(net1358),
    .A1(\vmem[479] ),
    .S(_06508_),
    .X(_01672_));
 or2_2 _22066_ (.A(net898),
    .B(_06413_),
    .X(_06509_));
 or4_1 _22067_ (.A(net783),
    .B(net622),
    .C(net871),
    .D(_06509_),
    .X(_06510_));
 mux2_1 _22068_ (.A0(net1368),
    .A1(\vmem[478] ),
    .S(_06510_),
    .X(_01673_));
 nand2_2 _22069_ (.A(net908),
    .B(_06416_),
    .Y(_06511_));
 or4_1 _22070_ (.A(net775),
    .B(net616),
    .C(net864),
    .D(_06511_),
    .X(_06512_));
 mux2_1 _22071_ (.A0(net1353),
    .A1(\vmem[477] ),
    .S(_06512_),
    .X(_01674_));
 or2_2 _22072_ (.A(net903),
    .B(_06419_),
    .X(_06513_));
 or4_1 _22073_ (.A(net796),
    .B(net635),
    .C(net882),
    .D(_06513_),
    .X(_06514_));
 mux2_1 _22074_ (.A0(net1386),
    .A1(\vmem[476] ),
    .S(_06514_),
    .X(_01675_));
 nand2_2 _22075_ (.A(net907),
    .B(_06422_),
    .Y(_06515_));
 or4_1 _22076_ (.A(net780),
    .B(net620),
    .C(net868),
    .D(_06515_),
    .X(_06516_));
 mux2_1 _22077_ (.A0(net1361),
    .A1(\vmem[475] ),
    .S(_06516_),
    .X(_01676_));
 or2_2 _22078_ (.A(net893),
    .B(_06425_),
    .X(_06517_));
 or4_1 _22079_ (.A(net771),
    .B(net614),
    .C(net862),
    .D(_06517_),
    .X(_06518_));
 mux2_1 _22080_ (.A0(net1346),
    .A1(\vmem[474] ),
    .S(_06518_),
    .X(_01677_));
 nand2_2 _22081_ (.A(net910),
    .B(_06428_),
    .Y(_06519_));
 or4_1 _22082_ (.A(net786),
    .B(net625),
    .C(net874),
    .D(_06519_),
    .X(_06520_));
 mux2_1 _22083_ (.A0(net1371),
    .A1(\vmem[473] ),
    .S(_06520_),
    .X(_01678_));
 nand2_2 _22084_ (.A(net906),
    .B(_06431_),
    .Y(_06521_));
 or4_1 _22085_ (.A(net763),
    .B(net610),
    .C(net857),
    .D(_06521_),
    .X(_06522_));
 mux2_1 _22086_ (.A0(net1336),
    .A1(\vmem[472] ),
    .S(_06522_),
    .X(_01679_));
 or2_2 _22087_ (.A(net895),
    .B(_06434_),
    .X(_06523_));
 or4_1 _22088_ (.A(net773),
    .B(net615),
    .C(net863),
    .D(_06523_),
    .X(_06524_));
 mux2_1 _22089_ (.A0(net1349),
    .A1(\vmem[471] ),
    .S(_06524_),
    .X(_01680_));
 or2_2 _22090_ (.A(net903),
    .B(_06437_),
    .X(_06525_));
 or4_1 _22091_ (.A(net797),
    .B(net636),
    .C(net883),
    .D(_06525_),
    .X(_06526_));
 mux2_1 _22092_ (.A0(net1390),
    .A1(\vmem[470] ),
    .S(_06526_),
    .X(_01681_));
 nand2_2 _22093_ (.A(net906),
    .B(_06440_),
    .Y(_06527_));
 or4_1 _22094_ (.A(net762),
    .B(net606),
    .C(net856),
    .D(_06527_),
    .X(_06528_));
 mux2_1 _22095_ (.A0(net1333),
    .A1(\vmem[469] ),
    .S(_06528_),
    .X(_01682_));
 or2_2 _22096_ (.A(net902),
    .B(_06443_),
    .X(_06529_));
 or4_1 _22097_ (.A(net793),
    .B(net631),
    .C(net880),
    .D(_06529_),
    .X(_06530_));
 mux2_1 _22098_ (.A0(net1380),
    .A1(\vmem[468] ),
    .S(_06530_),
    .X(_01683_));
 nand2_2 _22099_ (.A(net906),
    .B(_06446_),
    .Y(_06531_));
 or4_1 _22100_ (.A(net760),
    .B(net605),
    .C(net853),
    .D(_06531_),
    .X(_06532_));
 mux2_1 _22101_ (.A0(net1330),
    .A1(\vmem[467] ),
    .S(_06532_),
    .X(_01684_));
 or2_2 _22102_ (.A(net900),
    .B(_06449_),
    .X(_06533_));
 or4_1 _22103_ (.A(net795),
    .B(net630),
    .C(net880),
    .D(_06533_),
    .X(_06534_));
 mux2_1 _22104_ (.A0(net1381),
    .A1(\vmem[466] ),
    .S(_06534_),
    .X(_01685_));
 nand2_2 _22105_ (.A(net910),
    .B(_06452_),
    .Y(_06535_));
 or4_1 _22106_ (.A(net790),
    .B(net628),
    .C(net877),
    .D(_06535_),
    .X(_06536_));
 mux2_1 _22107_ (.A0(net1377),
    .A1(\vmem[465] ),
    .S(_06536_),
    .X(_01686_));
 nand2_2 _22108_ (.A(net906),
    .B(_06456_),
    .Y(_06537_));
 or4_1 _22109_ (.A(net766),
    .B(net612),
    .C(net859),
    .D(_06537_),
    .X(_06538_));
 mux2_1 _22110_ (.A0(net1341),
    .A1(\vmem[464] ),
    .S(_06538_),
    .X(_01687_));
 or2_2 _22111_ (.A(net896),
    .B(_06459_),
    .X(_06539_));
 or4_1 _22112_ (.A(net778),
    .B(net618),
    .C(net867),
    .D(_06539_),
    .X(_06540_));
 mux2_1 _22113_ (.A0(net1358),
    .A1(\vmem[463] ),
    .S(_06540_),
    .X(_01688_));
 or2_2 _22114_ (.A(net898),
    .B(_06462_),
    .X(_06541_));
 or4_1 _22115_ (.A(net783),
    .B(net622),
    .C(net870),
    .D(_06541_),
    .X(_06542_));
 mux2_1 _22116_ (.A0(net1368),
    .A1(\vmem[462] ),
    .S(_06542_),
    .X(_01689_));
 nand2_2 _22117_ (.A(net907),
    .B(_06465_),
    .Y(_06543_));
 or4_1 _22118_ (.A(net774),
    .B(net616),
    .C(net864),
    .D(_06543_),
    .X(_06544_));
 mux2_1 _22119_ (.A0(net1353),
    .A1(\vmem[461] ),
    .S(_06544_),
    .X(_01690_));
 or2_2 _22120_ (.A(net903),
    .B(_06468_),
    .X(_06545_));
 or4_1 _22121_ (.A(net796),
    .B(net635),
    .C(net882),
    .D(_06545_),
    .X(_06546_));
 mux2_1 _22122_ (.A0(net1386),
    .A1(\vmem[460] ),
    .S(_06546_),
    .X(_01691_));
 nand2_2 _22123_ (.A(net907),
    .B(_06471_),
    .Y(_06547_));
 or4_1 _22124_ (.A(net780),
    .B(net620),
    .C(net868),
    .D(_06547_),
    .X(_06548_));
 mux2_1 _22125_ (.A0(net1361),
    .A1(\vmem[459] ),
    .S(_06548_),
    .X(_01692_));
 or2_2 _22126_ (.A(net893),
    .B(_06474_),
    .X(_06549_));
 or4_1 _22127_ (.A(net770),
    .B(net614),
    .C(net862),
    .D(_06549_),
    .X(_06550_));
 mux2_1 _22128_ (.A0(net1345),
    .A1(\vmem[458] ),
    .S(_06550_),
    .X(_01693_));
 nand2_2 _22129_ (.A(net910),
    .B(_06477_),
    .Y(_06551_));
 or4_1 _22130_ (.A(net787),
    .B(net626),
    .C(net874),
    .D(_06551_),
    .X(_06552_));
 mux2_1 _22131_ (.A0(net1373),
    .A1(\vmem[457] ),
    .S(_06552_),
    .X(_01694_));
 nand2_2 _22132_ (.A(net906),
    .B(_06480_),
    .Y(_06553_));
 or4_1 _22133_ (.A(net764),
    .B(net610),
    .C(net855),
    .D(_06553_),
    .X(_06554_));
 mux2_1 _22134_ (.A0(net1336),
    .A1(\vmem[456] ),
    .S(_06554_),
    .X(_01695_));
 or2_2 _22135_ (.A(net895),
    .B(_06483_),
    .X(_06555_));
 or4_1 _22136_ (.A(net773),
    .B(net615),
    .C(net863),
    .D(_06555_),
    .X(_06556_));
 mux2_1 _22137_ (.A0(net1349),
    .A1(\vmem[455] ),
    .S(_06556_),
    .X(_01696_));
 or2_2 _22138_ (.A(net903),
    .B(_06486_),
    .X(_06557_));
 or4_1 _22139_ (.A(net797),
    .B(net636),
    .C(net883),
    .D(_06557_),
    .X(_06558_));
 mux2_1 _22140_ (.A0(net1392),
    .A1(\vmem[454] ),
    .S(_06558_),
    .X(_01697_));
 nand2_2 _22141_ (.A(net906),
    .B(_06489_),
    .Y(_06559_));
 or4_1 _22142_ (.A(net762),
    .B(net606),
    .C(net856),
    .D(_06559_),
    .X(_06560_));
 mux2_1 _22143_ (.A0(net1333),
    .A1(\vmem[453] ),
    .S(_06560_),
    .X(_01698_));
 or2_2 _22144_ (.A(net902),
    .B(_06492_),
    .X(_06561_));
 or4_1 _22145_ (.A(net793),
    .B(net631),
    .C(net879),
    .D(_06561_),
    .X(_06562_));
 mux2_1 _22146_ (.A0(net1383),
    .A1(\vmem[452] ),
    .S(_06562_),
    .X(_01699_));
 nand2_2 _22147_ (.A(net906),
    .B(_06495_),
    .Y(_06563_));
 or4_1 _22148_ (.A(net758),
    .B(net604),
    .C(net853),
    .D(_06563_),
    .X(_06564_));
 mux2_1 _22149_ (.A0(net1328),
    .A1(\vmem[451] ),
    .S(_06564_),
    .X(_01700_));
 or2_2 _22150_ (.A(net900),
    .B(_06498_),
    .X(_06565_));
 or4_1 _22151_ (.A(net792),
    .B(net630),
    .C(net880),
    .D(_06565_),
    .X(_06566_));
 mux2_1 _22152_ (.A0(net1381),
    .A1(\vmem[450] ),
    .S(_06566_),
    .X(_01701_));
 nand2_2 _22153_ (.A(net910),
    .B(_06501_),
    .Y(_06567_));
 or4_1 _22154_ (.A(net790),
    .B(net627),
    .C(net877),
    .D(_06567_),
    .X(_06568_));
 mux2_1 _22155_ (.A0(net1377),
    .A1(\vmem[449] ),
    .S(_06568_),
    .X(_01702_));
 nand2_2 _22156_ (.A(_03759_),
    .B(_06504_),
    .Y(_06569_));
 or4_1 _22157_ (.A(net766),
    .B(net612),
    .C(net860),
    .D(_06569_),
    .X(_06570_));
 mux2_1 _22158_ (.A0(net1341),
    .A1(\vmem[448] ),
    .S(_06570_),
    .X(_01703_));
 or4_1 _22159_ (.A(net736),
    .B(net619),
    .C(_06410_),
    .D(net867),
    .X(_06571_));
 mux2_1 _22160_ (.A0(net1359),
    .A1(\vmem[447] ),
    .S(_06571_),
    .X(_01704_));
 or4_1 _22161_ (.A(net740),
    .B(net623),
    .C(net871),
    .D(_06414_),
    .X(_06572_));
 mux2_1 _22162_ (.A0(net1368),
    .A1(\vmem[446] ),
    .S(_06572_),
    .X(_01705_));
 or4_1 _22163_ (.A(net739),
    .B(net621),
    .C(net865),
    .D(_06417_),
    .X(_06573_));
 mux2_1 _22164_ (.A0(net1365),
    .A1(\vmem[445] ),
    .S(_06573_),
    .X(_01706_));
 or4_1 _22165_ (.A(net753),
    .B(net634),
    .C(net882),
    .D(_06420_),
    .X(_06574_));
 mux2_1 _22166_ (.A0(net1386),
    .A1(\vmem[444] ),
    .S(_06574_),
    .X(_01707_));
 or4_1 _22167_ (.A(net738),
    .B(net624),
    .C(net869),
    .D(_06423_),
    .X(_06575_));
 mux2_1 _22168_ (.A0(net1362),
    .A1(\vmem[443] ),
    .S(_06575_),
    .X(_01708_));
 or4_1 _22169_ (.A(net725),
    .B(net611),
    .C(net858),
    .D(_06426_),
    .X(_06576_));
 mux2_1 _22170_ (.A0(net1339),
    .A1(\vmem[442] ),
    .S(_06576_),
    .X(_01709_));
 or4_1 _22171_ (.A(net743),
    .B(net625),
    .C(net876),
    .D(_06429_),
    .X(_06577_));
 mux2_1 _22172_ (.A0(net1372),
    .A1(\vmem[441] ),
    .S(_06577_),
    .X(_01710_));
 or4_1 _22173_ (.A(net724),
    .B(net610),
    .C(net858),
    .D(_06432_),
    .X(_06578_));
 mux2_1 _22174_ (.A0(net1337),
    .A1(\vmem[440] ),
    .S(_06578_),
    .X(_01711_));
 or4_1 _22175_ (.A(net734),
    .B(net616),
    .C(net864),
    .D(_06435_),
    .X(_06579_));
 mux2_1 _22176_ (.A0(net1352),
    .A1(\vmem[439] ),
    .S(_06579_),
    .X(_01712_));
 or4_1 _22177_ (.A(net755),
    .B(net636),
    .C(net883),
    .D(_06438_),
    .X(_06580_));
 mux2_1 _22178_ (.A0(net1390),
    .A1(\vmem[438] ),
    .S(_06580_),
    .X(_01713_));
 or4_1 _22179_ (.A(net723),
    .B(net606),
    .C(net856),
    .D(_06441_),
    .X(_06581_));
 mux2_1 _22180_ (.A0(net1333),
    .A1(\vmem[437] ),
    .S(_06581_),
    .X(_01714_));
 or4_1 _22181_ (.A(net749),
    .B(net630),
    .C(net880),
    .D(_06444_),
    .X(_06582_));
 mux2_1 _22182_ (.A0(net1380),
    .A1(\vmem[436] ),
    .S(_06582_),
    .X(_01715_));
 or4_1 _22183_ (.A(net721),
    .B(net605),
    .C(net855),
    .D(_06447_),
    .X(_06583_));
 mux2_1 _22184_ (.A0(net1330),
    .A1(\vmem[435] ),
    .S(_06583_),
    .X(_01716_));
 or4_1 _22185_ (.A(net749),
    .B(net633),
    .C(net875),
    .D(_06450_),
    .X(_06584_));
 mux2_1 _22186_ (.A0(net1381),
    .A1(\vmem[434] ),
    .S(_06584_),
    .X(_01717_));
 or4_1 _22187_ (.A(net747),
    .B(net628),
    .C(net878),
    .D(_06453_),
    .X(_06585_));
 mux2_1 _22188_ (.A0(net1377),
    .A1(\vmem[433] ),
    .S(_06585_),
    .X(_01718_));
 or4_1 _22189_ (.A(net728),
    .B(net612),
    .C(net859),
    .D(_06457_),
    .X(_06586_));
 mux2_1 _22190_ (.A0(net1343),
    .A1(\vmem[432] ),
    .S(_06586_),
    .X(_01719_));
 or4_1 _22191_ (.A(net735),
    .B(net619),
    .C(net866),
    .D(_06460_),
    .X(_06587_));
 mux2_1 _22192_ (.A0(net1357),
    .A1(\vmem[431] ),
    .S(_06587_),
    .X(_01720_));
 or4_1 _22193_ (.A(net740),
    .B(net622),
    .C(net870),
    .D(_06463_),
    .X(_06588_));
 mux2_1 _22194_ (.A0(net1369),
    .A1(\vmem[430] ),
    .S(_06588_),
    .X(_01721_));
 or4_1 _22195_ (.A(net739),
    .B(net621),
    .C(net872),
    .D(_06466_),
    .X(_06589_));
 mux2_1 _22196_ (.A0(net1365),
    .A1(\vmem[429] ),
    .S(_06589_),
    .X(_01722_));
 or4_1 _22197_ (.A(net753),
    .B(net634),
    .C(net882),
    .D(_06469_),
    .X(_06590_));
 mux2_1 _22198_ (.A0(net1386),
    .A1(\vmem[428] ),
    .S(_06590_),
    .X(_01723_));
 or4_1 _22199_ (.A(net738),
    .B(net620),
    .C(net869),
    .D(_06472_),
    .X(_06591_));
 mux2_1 _22200_ (.A0(net1362),
    .A1(\vmem[427] ),
    .S(_06591_),
    .X(_01724_));
 or4_1 _22201_ (.A(net726),
    .B(net611),
    .C(net858),
    .D(_06475_),
    .X(_06592_));
 mux2_1 _22202_ (.A0(net1339),
    .A1(\vmem[426] ),
    .S(_06592_),
    .X(_01725_));
 or4_1 _22203_ (.A(net745),
    .B(net625),
    .C(net876),
    .D(_06478_),
    .X(_06593_));
 mux2_1 _22204_ (.A0(net1393),
    .A1(\vmem[425] ),
    .S(_06593_),
    .X(_01726_));
 or4_1 _22205_ (.A(net724),
    .B(net610),
    .C(net857),
    .D(_06481_),
    .X(_06594_));
 mux2_1 _22206_ (.A0(net1337),
    .A1(\vmem[424] ),
    .S(_06594_),
    .X(_01727_));
 or4_1 _22207_ (.A(net734),
    .B(net616),
    .C(net864),
    .D(_06484_),
    .X(_06595_));
 mux2_1 _22208_ (.A0(net1352),
    .A1(\vmem[423] ),
    .S(_06595_),
    .X(_01728_));
 or4_1 _22209_ (.A(net754),
    .B(net637),
    .C(net883),
    .D(_06487_),
    .X(_06596_));
 mux2_1 _22210_ (.A0(net1392),
    .A1(\vmem[422] ),
    .S(_06596_),
    .X(_01729_));
 or4_1 _22211_ (.A(net723),
    .B(net606),
    .C(net856),
    .D(_06490_),
    .X(_06597_));
 mux2_1 _22212_ (.A0(net1333),
    .A1(\vmem[421] ),
    .S(_06597_),
    .X(_01730_));
 or4_1 _22213_ (.A(net752),
    .B(net630),
    .C(net880),
    .D(_06493_),
    .X(_06598_));
 mux2_1 _22214_ (.A0(net1381),
    .A1(\vmem[420] ),
    .S(_06598_),
    .X(_01731_));
 or4_1 _22215_ (.A(net721),
    .B(net605),
    .C(net853),
    .D(_06496_),
    .X(_06599_));
 mux2_1 _22216_ (.A0(net1330),
    .A1(\vmem[419] ),
    .S(_06599_),
    .X(_01732_));
 or4_1 _22217_ (.A(net752),
    .B(net630),
    .C(net875),
    .D(_06499_),
    .X(_06600_));
 mux2_1 _22218_ (.A0(net1381),
    .A1(\vmem[418] ),
    .S(_06600_),
    .X(_01733_));
 or4_1 _22219_ (.A(net747),
    .B(net628),
    .C(net878),
    .D(_06502_),
    .X(_06601_));
 mux2_1 _22220_ (.A0(net1377),
    .A1(\vmem[417] ),
    .S(_06601_),
    .X(_01734_));
 or4_1 _22221_ (.A(net728),
    .B(net612),
    .C(net859),
    .D(_06505_),
    .X(_06602_));
 mux2_1 _22222_ (.A0(net1343),
    .A1(\vmem[416] ),
    .S(_06602_),
    .X(_01735_));
 or4_1 _22223_ (.A(net735),
    .B(net618),
    .C(net867),
    .D(_06507_),
    .X(_06603_));
 mux2_1 _22224_ (.A0(net1359),
    .A1(\vmem[415] ),
    .S(_06603_),
    .X(_01736_));
 or4_1 _22225_ (.A(net741),
    .B(net622),
    .C(net871),
    .D(_06509_),
    .X(_06604_));
 mux2_1 _22226_ (.A0(net1369),
    .A1(\vmem[414] ),
    .S(_06604_),
    .X(_01737_));
 or4_1 _22227_ (.A(net733),
    .B(net616),
    .C(net864),
    .D(_06511_),
    .X(_06605_));
 mux2_1 _22228_ (.A0(net1353),
    .A1(\vmem[413] ),
    .S(_06605_),
    .X(_01738_));
 or4_1 _22229_ (.A(net753),
    .B(net634),
    .C(net882),
    .D(_06513_),
    .X(_06606_));
 mux2_1 _22230_ (.A0(net1389),
    .A1(\vmem[412] ),
    .S(_06606_),
    .X(_01739_));
 or4_1 _22231_ (.A(net738),
    .B(net620),
    .C(net869),
    .D(_06515_),
    .X(_06607_));
 mux2_1 _22232_ (.A0(net1361),
    .A1(\vmem[411] ),
    .S(_06607_),
    .X(_01740_));
 or4_1 _22233_ (.A(net730),
    .B(net614),
    .C(net861),
    .D(_06517_),
    .X(_06608_));
 mux2_1 _22234_ (.A0(net1345),
    .A1(\vmem[410] ),
    .S(_06608_),
    .X(_01741_));
 or4_1 _22235_ (.A(net743),
    .B(net625),
    .C(net874),
    .D(_06519_),
    .X(_06609_));
 mux2_1 _22236_ (.A0(net1371),
    .A1(\vmem[409] ),
    .S(_06609_),
    .X(_01742_));
 or4_1 _22237_ (.A(net724),
    .B(net609),
    .C(net857),
    .D(_06521_),
    .X(_06610_));
 mux2_1 _22238_ (.A0(net1335),
    .A1(\vmem[408] ),
    .S(_06610_),
    .X(_01743_));
 or4_1 _22239_ (.A(net731),
    .B(net615),
    .C(net863),
    .D(_06523_),
    .X(_06611_));
 mux2_1 _22240_ (.A0(net1350),
    .A1(\vmem[407] ),
    .S(_06611_),
    .X(_01744_));
 or4_1 _22241_ (.A(net755),
    .B(net636),
    .C(net883),
    .D(_06525_),
    .X(_06612_));
 mux2_1 _22242_ (.A0(net1390),
    .A1(\vmem[406] ),
    .S(_06612_),
    .X(_01745_));
 or4_1 _22243_ (.A(net723),
    .B(net606),
    .C(net856),
    .D(_06527_),
    .X(_06613_));
 mux2_1 _22244_ (.A0(net1333),
    .A1(\vmem[405] ),
    .S(_06613_),
    .X(_01746_));
 or4_1 _22245_ (.A(net750),
    .B(net631),
    .C(net879),
    .D(_06529_),
    .X(_06614_));
 mux2_1 _22246_ (.A0(net1383),
    .A1(\vmem[404] ),
    .S(_06614_),
    .X(_01747_));
 or4_1 _22247_ (.A(net721),
    .B(net605),
    .C(net853),
    .D(_06531_),
    .X(_06615_));
 mux2_1 _22248_ (.A0(net1332),
    .A1(\vmem[403] ),
    .S(_06615_),
    .X(_01748_));
 or4_1 _22249_ (.A(net749),
    .B(net630),
    .C(net880),
    .D(_06533_),
    .X(_06616_));
 mux2_1 _22250_ (.A0(net1382),
    .A1(\vmem[402] ),
    .S(_06616_),
    .X(_01749_));
 or4_1 _22251_ (.A(net747),
    .B(net628),
    .C(net878),
    .D(_06535_),
    .X(_06617_));
 mux2_1 _22252_ (.A0(net1377),
    .A1(\vmem[401] ),
    .S(_06617_),
    .X(_01750_));
 or4_1 _22253_ (.A(net727),
    .B(net612),
    .C(net860),
    .D(_06537_),
    .X(_06618_));
 mux2_1 _22254_ (.A0(net1341),
    .A1(\vmem[400] ),
    .S(_06618_),
    .X(_01751_));
 or4_1 _22255_ (.A(net736),
    .B(net618),
    .C(net867),
    .D(_06539_),
    .X(_06619_));
 mux2_1 _22256_ (.A0(net1358),
    .A1(\vmem[399] ),
    .S(_06619_),
    .X(_01752_));
 or4_1 _22257_ (.A(net740),
    .B(net622),
    .C(net871),
    .D(_06541_),
    .X(_06620_));
 mux2_1 _22258_ (.A0(net1369),
    .A1(\vmem[398] ),
    .S(_06620_),
    .X(_01753_));
 or4_1 _22259_ (.A(net734),
    .B(net617),
    .C(net864),
    .D(_06543_),
    .X(_06621_));
 mux2_1 _22260_ (.A0(net1353),
    .A1(\vmem[397] ),
    .S(_06621_),
    .X(_01754_));
 or4_1 _22261_ (.A(net753),
    .B(net635),
    .C(net882),
    .D(_06545_),
    .X(_06622_));
 mux2_1 _22262_ (.A0(net1386),
    .A1(\vmem[396] ),
    .S(_06622_),
    .X(_01755_));
 or4_1 _22263_ (.A(net738),
    .B(net620),
    .C(net869),
    .D(_06547_),
    .X(_06623_));
 mux2_1 _22264_ (.A0(net1362),
    .A1(\vmem[395] ),
    .S(_06623_),
    .X(_01756_));
 or4_1 _22265_ (.A(net730),
    .B(net614),
    .C(net861),
    .D(_06549_),
    .X(_06624_));
 mux2_1 _22266_ (.A0(net1345),
    .A1(\vmem[394] ),
    .S(_06624_),
    .X(_01757_));
 or4_1 _22267_ (.A(net743),
    .B(net625),
    .C(net874),
    .D(_06551_),
    .X(_06625_));
 mux2_1 _22268_ (.A0(net1372),
    .A1(\vmem[393] ),
    .S(_06625_),
    .X(_01758_));
 or4_1 _22269_ (.A(net724),
    .B(net610),
    .C(net857),
    .D(_06553_),
    .X(_06626_));
 mux2_1 _22270_ (.A0(net1337),
    .A1(\vmem[392] ),
    .S(_06626_),
    .X(_01759_));
 or4_1 _22271_ (.A(net731),
    .B(net615),
    .C(net863),
    .D(_06555_),
    .X(_06627_));
 mux2_1 _22272_ (.A0(net1349),
    .A1(\vmem[391] ),
    .S(_06627_),
    .X(_01760_));
 or4_1 _22273_ (.A(net755),
    .B(net636),
    .C(net883),
    .D(_06557_),
    .X(_06628_));
 mux2_1 _22274_ (.A0(net1390),
    .A1(\vmem[390] ),
    .S(_06628_),
    .X(_01761_));
 or4_1 _22275_ (.A(net723),
    .B(net606),
    .C(net856),
    .D(_06559_),
    .X(_06629_));
 mux2_1 _22276_ (.A0(net1333),
    .A1(\vmem[389] ),
    .S(_06629_),
    .X(_01762_));
 or4_1 _22277_ (.A(net750),
    .B(net632),
    .C(net879),
    .D(_06561_),
    .X(_06630_));
 mux2_1 _22278_ (.A0(net1383),
    .A1(\vmem[388] ),
    .S(_06630_),
    .X(_01763_));
 or4_1 _22279_ (.A(net721),
    .B(net605),
    .C(net854),
    .D(_06563_),
    .X(_06631_));
 mux2_1 _22280_ (.A0(net1330),
    .A1(\vmem[387] ),
    .S(_06631_),
    .X(_01764_));
 or4_1 _22281_ (.A(net749),
    .B(net630),
    .C(net880),
    .D(_06565_),
    .X(_06632_));
 mux2_1 _22282_ (.A0(net1381),
    .A1(\vmem[386] ),
    .S(_06632_),
    .X(_01765_));
 or4_1 _22283_ (.A(net746),
    .B(net627),
    .C(net877),
    .D(_06567_),
    .X(_06633_));
 mux2_1 _22284_ (.A0(net1376),
    .A1(\vmem[385] ),
    .S(_06633_),
    .X(_01766_));
 or4_1 _22285_ (.A(net727),
    .B(net612),
    .C(net860),
    .D(_06569_),
    .X(_06634_));
 mux2_1 _22286_ (.A0(net1341),
    .A1(\vmem[384] ),
    .S(_06634_),
    .X(_01767_));
 or4_1 _22287_ (.A(net777),
    .B(net655),
    .C(_06410_),
    .D(net866),
    .X(_06635_));
 mux2_1 _22288_ (.A0(net1356),
    .A1(\vmem[383] ),
    .S(_06635_),
    .X(_01768_));
 or4_1 _22289_ (.A(net783),
    .B(net659),
    .C(net870),
    .D(_06414_),
    .X(_06636_));
 mux2_1 _22290_ (.A0(net1367),
    .A1(\vmem[382] ),
    .S(_06636_),
    .X(_01769_));
 or4_1 _22291_ (.A(net781),
    .B(net661),
    .C(net872),
    .D(_06417_),
    .X(_06637_));
 mux2_1 _22292_ (.A0(net1364),
    .A1(\vmem[381] ),
    .S(_06637_),
    .X(_01770_));
 or4_1 _22293_ (.A(net796),
    .B(net671),
    .C(net881),
    .D(_06420_),
    .X(_06638_));
 mux2_1 _22294_ (.A0(net1387),
    .A1(\vmem[380] ),
    .S(_06638_),
    .X(_01771_));
 or4_1 _22295_ (.A(net779),
    .B(net658),
    .C(net868),
    .D(_06423_),
    .X(_06639_));
 mux2_1 _22296_ (.A0(net1360),
    .A1(\vmem[379] ),
    .S(_06639_),
    .X(_01772_));
 or4_1 _22297_ (.A(net770),
    .B(net650),
    .C(net862),
    .D(_06426_),
    .X(_06640_));
 mux2_1 _22298_ (.A0(net1347),
    .A1(\vmem[378] ),
    .S(_06640_),
    .X(_01773_));
 or4_1 _22299_ (.A(net786),
    .B(net664),
    .C(net874),
    .D(_06429_),
    .X(_06641_));
 mux2_1 _22300_ (.A0(net1372),
    .A1(\vmem[377] ),
    .S(_06641_),
    .X(_01774_));
 or4_1 _22301_ (.A(net768),
    .B(net644),
    .C(net858),
    .D(_06432_),
    .X(_06642_));
 mux2_1 _22302_ (.A0(net1339),
    .A1(\vmem[376] ),
    .S(_06642_),
    .X(_01775_));
 or4_1 _22303_ (.A(net774),
    .B(net652),
    .C(net865),
    .D(_06435_),
    .X(_06643_));
 mux2_1 _22304_ (.A0(net1352),
    .A1(\vmem[375] ),
    .S(_06643_),
    .X(_01776_));
 or4_1 _22305_ (.A(net797),
    .B(net672),
    .C(net884),
    .D(_06438_),
    .X(_06644_));
 mux2_1 _22306_ (.A0(net1391),
    .A1(\vmem[374] ),
    .S(_06644_),
    .X(_01777_));
 or4_1 _22307_ (.A(net760),
    .B(net642),
    .C(net855),
    .D(_06441_),
    .X(_06645_));
 mux2_1 _22308_ (.A0(net1331),
    .A1(\vmem[373] ),
    .S(_06645_),
    .X(_01778_));
 or4_1 _22309_ (.A(net794),
    .B(net668),
    .C(net879),
    .D(_06444_),
    .X(_06646_));
 mux2_1 _22310_ (.A0(net1385),
    .A1(\vmem[372] ),
    .S(_06646_),
    .X(_01779_));
 or4_1 _22311_ (.A(net759),
    .B(net640),
    .C(net853),
    .D(_06447_),
    .X(_06647_));
 mux2_1 _22312_ (.A0(net1328),
    .A1(\vmem[371] ),
    .S(_06647_),
    .X(_01780_));
 or4_1 _22313_ (.A(net787),
    .B(net663),
    .C(net875),
    .D(_06450_),
    .X(_06648_));
 mux2_1 _22314_ (.A0(net1373),
    .A1(\vmem[370] ),
    .S(_06648_),
    .X(_01781_));
 or4_1 _22315_ (.A(net788),
    .B(net663),
    .C(net875),
    .D(_06453_),
    .X(_06649_));
 mux2_1 _22316_ (.A0(net1374),
    .A1(\vmem[369] ),
    .S(_06649_),
    .X(_01782_));
 or4_1 _22317_ (.A(net767),
    .B(net646),
    .C(net859),
    .D(_06457_),
    .X(_06650_));
 mux2_1 _22318_ (.A0(net1342),
    .A1(\vmem[368] ),
    .S(_06650_),
    .X(_01783_));
 or4_1 _22319_ (.A(net777),
    .B(net655),
    .C(net866),
    .D(_06460_),
    .X(_06651_));
 mux2_1 _22320_ (.A0(net1356),
    .A1(\vmem[367] ),
    .S(_06651_),
    .X(_01784_));
 or4_1 _22321_ (.A(net782),
    .B(net659),
    .C(net870),
    .D(_06463_),
    .X(_06652_));
 mux2_1 _22322_ (.A0(net1367),
    .A1(\vmem[366] ),
    .S(_06652_),
    .X(_01785_));
 or4_1 _22323_ (.A(net781),
    .B(net661),
    .C(net872),
    .D(_06466_),
    .X(_06653_));
 mux2_1 _22324_ (.A0(net1364),
    .A1(\vmem[365] ),
    .S(_06653_),
    .X(_01786_));
 or4_1 _22325_ (.A(net796),
    .B(net671),
    .C(net881),
    .D(_06469_),
    .X(_06654_));
 mux2_1 _22326_ (.A0(net1387),
    .A1(\vmem[364] ),
    .S(_06654_),
    .X(_01787_));
 or4_1 _22327_ (.A(net780),
    .B(net658),
    .C(net869),
    .D(_06472_),
    .X(_06655_));
 mux2_1 _22328_ (.A0(net1361),
    .A1(\vmem[363] ),
    .S(_06655_),
    .X(_01788_));
 or4_1 _22329_ (.A(net770),
    .B(net650),
    .C(net862),
    .D(_06475_),
    .X(_06656_));
 mux2_1 _22330_ (.A0(net1347),
    .A1(\vmem[362] ),
    .S(_06656_),
    .X(_01789_));
 or4_1 _22331_ (.A(net786),
    .B(net664),
    .C(net874),
    .D(_06478_),
    .X(_06657_));
 mux2_1 _22332_ (.A0(net1371),
    .A1(\vmem[361] ),
    .S(_06657_),
    .X(_01790_));
 or4_1 _22333_ (.A(net768),
    .B(net647),
    .C(net857),
    .D(_06481_),
    .X(_06658_));
 mux2_1 _22334_ (.A0(net1339),
    .A1(\vmem[360] ),
    .S(_06658_),
    .X(_01791_));
 or4_1 _22335_ (.A(net774),
    .B(net652),
    .C(net865),
    .D(_06484_),
    .X(_06659_));
 mux2_1 _22336_ (.A0(net1352),
    .A1(\vmem[359] ),
    .S(_06659_),
    .X(_01792_));
 or4_1 _22337_ (.A(net797),
    .B(net672),
    .C(net884),
    .D(_06487_),
    .X(_06660_));
 mux2_1 _22338_ (.A0(net1391),
    .A1(\vmem[358] ),
    .S(_06660_),
    .X(_01793_));
 or4_1 _22339_ (.A(net760),
    .B(net642),
    .C(net854),
    .D(_06490_),
    .X(_06661_));
 mux2_1 _22340_ (.A0(net1331),
    .A1(\vmem[357] ),
    .S(_06661_),
    .X(_01794_));
 or4_1 _22341_ (.A(net794),
    .B(net668),
    .C(net879),
    .D(_06493_),
    .X(_06662_));
 mux2_1 _22342_ (.A0(net1385),
    .A1(\vmem[356] ),
    .S(_06662_),
    .X(_01795_));
 or4_1 _22343_ (.A(net760),
    .B(net641),
    .C(net853),
    .D(_06496_),
    .X(_06663_));
 mux2_1 _22344_ (.A0(net1330),
    .A1(\vmem[355] ),
    .S(_06663_),
    .X(_01796_));
 or4_1 _22345_ (.A(net788),
    .B(net663),
    .C(net875),
    .D(_06499_),
    .X(_06664_));
 mux2_1 _22346_ (.A0(net1374),
    .A1(\vmem[354] ),
    .S(_06664_),
    .X(_01797_));
 or4_1 _22347_ (.A(net789),
    .B(net666),
    .C(net878),
    .D(_06502_),
    .X(_06665_));
 mux2_1 _22348_ (.A0(net1374),
    .A1(\vmem[353] ),
    .S(_06665_),
    .X(_01798_));
 or4_1 _22349_ (.A(net767),
    .B(net646),
    .C(net859),
    .D(_06505_),
    .X(_06666_));
 mux2_1 _22350_ (.A0(net1342),
    .A1(\vmem[352] ),
    .S(_06666_),
    .X(_01799_));
 or4_1 _22351_ (.A(net777),
    .B(net656),
    .C(net866),
    .D(_06507_),
    .X(_06667_));
 mux2_1 _22352_ (.A0(net1356),
    .A1(\vmem[351] ),
    .S(_06667_),
    .X(_01800_));
 or4_1 _22353_ (.A(net782),
    .B(net660),
    .C(net870),
    .D(_06509_),
    .X(_06668_));
 mux2_1 _22354_ (.A0(net1369),
    .A1(\vmem[350] ),
    .S(_06668_),
    .X(_01801_));
 or4_1 _22355_ (.A(net781),
    .B(net661),
    .C(net872),
    .D(_06511_),
    .X(_06669_));
 mux2_1 _22356_ (.A0(net1364),
    .A1(\vmem[349] ),
    .S(_06669_),
    .X(_01802_));
 or4_1 _22357_ (.A(net799),
    .B(net674),
    .C(net881),
    .D(_06513_),
    .X(_06670_));
 mux2_1 _22358_ (.A0(net1388),
    .A1(\vmem[348] ),
    .S(_06670_),
    .X(_01803_));
 or4_1 _22359_ (.A(net780),
    .B(net658),
    .C(net869),
    .D(_06515_),
    .X(_06671_));
 mux2_1 _22360_ (.A0(net1361),
    .A1(\vmem[347] ),
    .S(_06671_),
    .X(_01804_));
 or4_1 _22361_ (.A(net772),
    .B(net650),
    .C(net863),
    .D(_06517_),
    .X(_06672_));
 mux2_1 _22362_ (.A0(net1347),
    .A1(\vmem[346] ),
    .S(_06672_),
    .X(_01805_));
 or4_1 _22363_ (.A(net775),
    .B(net652),
    .C(net865),
    .D(_06519_),
    .X(_06673_));
 mux2_1 _22364_ (.A0(net1351),
    .A1(\vmem[345] ),
    .S(_06673_),
    .X(_01806_));
 or4_1 _22365_ (.A(net765),
    .B(net643),
    .C(net858),
    .D(_06521_),
    .X(_06674_));
 mux2_1 _22366_ (.A0(net1338),
    .A1(\vmem[344] ),
    .S(_06674_),
    .X(_01807_));
 or4_1 _22367_ (.A(net772),
    .B(net651),
    .C(net862),
    .D(_06523_),
    .X(_06675_));
 mux2_1 _22368_ (.A0(net1349),
    .A1(\vmem[343] ),
    .S(_06675_),
    .X(_01808_));
 or4_1 _22369_ (.A(net798),
    .B(net672),
    .C(net882),
    .D(_06525_),
    .X(_06676_));
 mux2_1 _22370_ (.A0(net1387),
    .A1(\vmem[342] ),
    .S(_06676_),
    .X(_01809_));
 or4_1 _22371_ (.A(net763),
    .B(net644),
    .C(net854),
    .D(_06527_),
    .X(_06677_));
 mux2_1 _22372_ (.A0(net1336),
    .A1(\vmem[341] ),
    .S(_06677_),
    .X(_01810_));
 or4_1 _22373_ (.A(net794),
    .B(net668),
    .C(net879),
    .D(_06529_),
    .X(_06678_));
 mux2_1 _22374_ (.A0(net1384),
    .A1(\vmem[340] ),
    .S(_06678_),
    .X(_01811_));
 or4_1 _22375_ (.A(net760),
    .B(net641),
    .C(net854),
    .D(_06531_),
    .X(_06679_));
 mux2_1 _22376_ (.A0(net1330),
    .A1(\vmem[339] ),
    .S(_06679_),
    .X(_01812_));
 or4_1 _22377_ (.A(net787),
    .B(net663),
    .C(net876),
    .D(_06533_),
    .X(_06680_));
 mux2_1 _22378_ (.A0(net1375),
    .A1(\vmem[338] ),
    .S(_06680_),
    .X(_01813_));
 or4_1 _22379_ (.A(net787),
    .B(net665),
    .C(net875),
    .D(_06535_),
    .X(_06681_));
 mux2_1 _22380_ (.A0(net1375),
    .A1(\vmem[337] ),
    .S(_06681_),
    .X(_01814_));
 or4_1 _22381_ (.A(net764),
    .B(net644),
    .C(net857),
    .D(_06537_),
    .X(_06682_));
 mux2_1 _22382_ (.A0(net1336),
    .A1(\vmem[336] ),
    .S(_06682_),
    .X(_01815_));
 or4_1 _22383_ (.A(net777),
    .B(net655),
    .C(net866),
    .D(_06539_),
    .X(_06683_));
 mux2_1 _22384_ (.A0(net1356),
    .A1(\vmem[335] ),
    .S(_06683_),
    .X(_01816_));
 or4_1 _22385_ (.A(net782),
    .B(net660),
    .C(net870),
    .D(_06541_),
    .X(_06684_));
 mux2_1 _22386_ (.A0(net1369),
    .A1(\vmem[334] ),
    .S(_06684_),
    .X(_01817_));
 or4_1 _22387_ (.A(net778),
    .B(net656),
    .C(net867),
    .D(_06543_),
    .X(_06685_));
 mux2_1 _22388_ (.A0(net1358),
    .A1(\vmem[333] ),
    .S(_06685_),
    .X(_01818_));
 or4_1 _22389_ (.A(net799),
    .B(net674),
    .C(net881),
    .D(_06545_),
    .X(_06686_));
 mux2_1 _22390_ (.A0(net1388),
    .A1(\vmem[332] ),
    .S(_06686_),
    .X(_01819_));
 or4_1 _22391_ (.A(net779),
    .B(net657),
    .C(net868),
    .D(_06547_),
    .X(_06687_));
 mux2_1 _22392_ (.A0(net1360),
    .A1(\vmem[331] ),
    .S(_06687_),
    .X(_01820_));
 or4_1 _22393_ (.A(net772),
    .B(net650),
    .C(net862),
    .D(_06549_),
    .X(_06688_));
 mux2_1 _22394_ (.A0(net1347),
    .A1(\vmem[330] ),
    .S(_06688_),
    .X(_01821_));
 or4_1 _22395_ (.A(net775),
    .B(net652),
    .C(net865),
    .D(_06551_),
    .X(_06689_));
 mux2_1 _22396_ (.A0(net1355),
    .A1(\vmem[329] ),
    .S(_06689_),
    .X(_01822_));
 or4_1 _22397_ (.A(net765),
    .B(net643),
    .C(net857),
    .D(_06553_),
    .X(_06690_));
 mux2_1 _22398_ (.A0(net1338),
    .A1(\vmem[328] ),
    .S(_06690_),
    .X(_01823_));
 or4_1 _22399_ (.A(net772),
    .B(net651),
    .C(net862),
    .D(_06555_),
    .X(_06691_));
 mux2_1 _22400_ (.A0(net1349),
    .A1(\vmem[327] ),
    .S(_06691_),
    .X(_01824_));
 or4_1 _22401_ (.A(net797),
    .B(net672),
    .C(net881),
    .D(_06557_),
    .X(_06692_));
 mux2_1 _22402_ (.A0(net1388),
    .A1(\vmem[326] ),
    .S(_06692_),
    .X(_01825_));
 or4_1 _22403_ (.A(net764),
    .B(net644),
    .C(net854),
    .D(_06559_),
    .X(_06693_));
 mux2_1 _22404_ (.A0(net1336),
    .A1(\vmem[325] ),
    .S(_06693_),
    .X(_01826_));
 or4_1 _22405_ (.A(net794),
    .B(net668),
    .C(net879),
    .D(_06561_),
    .X(_06694_));
 mux2_1 _22406_ (.A0(net1384),
    .A1(\vmem[324] ),
    .S(_06694_),
    .X(_01827_));
 or4_1 _22407_ (.A(net760),
    .B(net641),
    .C(net854),
    .D(_06563_),
    .X(_06695_));
 mux2_1 _22408_ (.A0(net1330),
    .A1(\vmem[323] ),
    .S(_06695_),
    .X(_01828_));
 or4_1 _22409_ (.A(net787),
    .B(net665),
    .C(net876),
    .D(_06565_),
    .X(_06696_));
 mux2_1 _22410_ (.A0(net1375),
    .A1(\vmem[322] ),
    .S(_06696_),
    .X(_01829_));
 or4_1 _22411_ (.A(net789),
    .B(net666),
    .C(net877),
    .D(_06567_),
    .X(_06697_));
 mux2_1 _22412_ (.A0(net1378),
    .A1(\vmem[321] ),
    .S(_06697_),
    .X(_01830_));
 or4_1 _22413_ (.A(net766),
    .B(net645),
    .C(net859),
    .D(_06569_),
    .X(_06698_));
 mux2_1 _22414_ (.A0(net1340),
    .A1(\vmem[320] ),
    .S(_06698_),
    .X(_01831_));
 or4_1 _22415_ (.A(net735),
    .B(net656),
    .C(_06410_),
    .D(net866),
    .X(_06699_));
 mux2_1 _22416_ (.A0(net1357),
    .A1(\vmem[319] ),
    .S(_06699_),
    .X(_01832_));
 or4_1 _22417_ (.A(net740),
    .B(net659),
    .C(net870),
    .D(_06414_),
    .X(_06700_));
 mux2_1 _22418_ (.A0(net1367),
    .A1(\vmem[318] ),
    .S(_06700_),
    .X(_01833_));
 or4_1 _22419_ (.A(net739),
    .B(net661),
    .C(net872),
    .D(_06417_),
    .X(_06701_));
 mux2_1 _22420_ (.A0(net1364),
    .A1(\vmem[317] ),
    .S(_06701_),
    .X(_01834_));
 or4_1 _22421_ (.A(net753),
    .B(net671),
    .C(net881),
    .D(_06420_),
    .X(_06702_));
 mux2_1 _22422_ (.A0(net1387),
    .A1(\vmem[316] ),
    .S(_06702_),
    .X(_01835_));
 or4_1 _22423_ (.A(net737),
    .B(net658),
    .C(net868),
    .D(_06423_),
    .X(_06703_));
 mux2_1 _22424_ (.A0(net1362),
    .A1(\vmem[315] ),
    .S(_06703_),
    .X(_01836_));
 or4_1 _22425_ (.A(net732),
    .B(net651),
    .C(net862),
    .D(_06426_),
    .X(_06704_));
 mux2_1 _22426_ (.A0(net1349),
    .A1(\vmem[314] ),
    .S(_06704_),
    .X(_01837_));
 or4_1 _22427_ (.A(net743),
    .B(net664),
    .C(net874),
    .D(_06429_),
    .X(_06705_));
 mux2_1 _22428_ (.A0(net1372),
    .A1(\vmem[313] ),
    .S(_06705_),
    .X(_01838_));
 or4_1 _22429_ (.A(net726),
    .B(net647),
    .C(net858),
    .D(_06432_),
    .X(_06706_));
 mux2_1 _22430_ (.A0(net1339),
    .A1(\vmem[312] ),
    .S(_06706_),
    .X(_01839_));
 or4_1 _22431_ (.A(net734),
    .B(net653),
    .C(net864),
    .D(_06435_),
    .X(_06707_));
 mux2_1 _22432_ (.A0(net1353),
    .A1(\vmem[311] ),
    .S(_06707_),
    .X(_01840_));
 or4_1 _22433_ (.A(net754),
    .B(net672),
    .C(net883),
    .D(_06438_),
    .X(_06708_));
 mux2_1 _22434_ (.A0(net1391),
    .A1(\vmem[310] ),
    .S(_06708_),
    .X(_01841_));
 or4_1 _22435_ (.A(net723),
    .B(net647),
    .C(net856),
    .D(_06441_),
    .X(_06709_));
 mux2_1 _22436_ (.A0(net1333),
    .A1(\vmem[309] ),
    .S(_06709_),
    .X(_01842_));
 or4_1 _22437_ (.A(net751),
    .B(net668),
    .C(net879),
    .D(_06444_),
    .X(_06710_));
 mux2_1 _22438_ (.A0(net1385),
    .A1(\vmem[308] ),
    .S(_06710_),
    .X(_01843_));
 or4_1 _22439_ (.A(net721),
    .B(net641),
    .C(net853),
    .D(_06447_),
    .X(_06711_));
 mux2_1 _22440_ (.A0(net1330),
    .A1(\vmem[307] ),
    .S(_06711_),
    .X(_01844_));
 or4_1 _22441_ (.A(net744),
    .B(net663),
    .C(net875),
    .D(_06450_),
    .X(_06712_));
 mux2_1 _22442_ (.A0(net1373),
    .A1(\vmem[306] ),
    .S(_06712_),
    .X(_01845_));
 or4_1 _22443_ (.A(net746),
    .B(net666),
    .C(net877),
    .D(_06453_),
    .X(_06713_));
 mux2_1 _22444_ (.A0(net1376),
    .A1(\vmem[305] ),
    .S(_06713_),
    .X(_01846_));
 or4_1 _22445_ (.A(net728),
    .B(net646),
    .C(net859),
    .D(_06457_),
    .X(_06714_));
 mux2_1 _22446_ (.A0(net1342),
    .A1(\vmem[304] ),
    .S(_06714_),
    .X(_01847_));
 or4_1 _22447_ (.A(net735),
    .B(net656),
    .C(net866),
    .D(_06460_),
    .X(_06715_));
 mux2_1 _22448_ (.A0(net1357),
    .A1(\vmem[303] ),
    .S(_06715_),
    .X(_01848_));
 or4_1 _22449_ (.A(net740),
    .B(net659),
    .C(net870),
    .D(_06463_),
    .X(_06716_));
 mux2_1 _22450_ (.A0(net1367),
    .A1(\vmem[302] ),
    .S(_06716_),
    .X(_01849_));
 or4_1 _22451_ (.A(net739),
    .B(net661),
    .C(net872),
    .D(_06466_),
    .X(_06717_));
 mux2_1 _22452_ (.A0(net1364),
    .A1(\vmem[301] ),
    .S(_06717_),
    .X(_01850_));
 or4_1 _22453_ (.A(net753),
    .B(net671),
    .C(net881),
    .D(_06469_),
    .X(_06718_));
 mux2_1 _22454_ (.A0(net1387),
    .A1(\vmem[300] ),
    .S(_06718_),
    .X(_01851_));
 or4_1 _22455_ (.A(net737),
    .B(net657),
    .C(net868),
    .D(_06472_),
    .X(_06719_));
 mux2_1 _22456_ (.A0(net1362),
    .A1(\vmem[299] ),
    .S(_06719_),
    .X(_01852_));
 or4_1 _22457_ (.A(net731),
    .B(net650),
    .C(net862),
    .D(_06475_),
    .X(_06720_));
 mux2_1 _22458_ (.A0(net1347),
    .A1(\vmem[298] ),
    .S(_06720_),
    .X(_01853_));
 or4_1 _22459_ (.A(net744),
    .B(net663),
    .C(net874),
    .D(_06478_),
    .X(_06721_));
 mux2_1 _22460_ (.A0(net1373),
    .A1(\vmem[297] ),
    .S(_06721_),
    .X(_01854_));
 or4_1 _22461_ (.A(net726),
    .B(net643),
    .C(net857),
    .D(_06481_),
    .X(_06722_));
 mux2_1 _22462_ (.A0(net1339),
    .A1(\vmem[296] ),
    .S(_06722_),
    .X(_01855_));
 or4_1 _22463_ (.A(net733),
    .B(net653),
    .C(net864),
    .D(_06484_),
    .X(_06723_));
 mux2_1 _22464_ (.A0(net1353),
    .A1(\vmem[295] ),
    .S(_06723_),
    .X(_01856_));
 or4_1 _22465_ (.A(net754),
    .B(net672),
    .C(net884),
    .D(_06487_),
    .X(_06724_));
 mux2_1 _22466_ (.A0(net1391),
    .A1(\vmem[294] ),
    .S(_06724_),
    .X(_01857_));
 or4_1 _22467_ (.A(net729),
    .B(net642),
    .C(net854),
    .D(_06490_),
    .X(_06725_));
 mux2_1 _22468_ (.A0(net1331),
    .A1(\vmem[293] ),
    .S(_06725_),
    .X(_01858_));
 or4_1 _22469_ (.A(net750),
    .B(net669),
    .C(net885),
    .D(_06493_),
    .X(_06726_));
 mux2_1 _22470_ (.A0(net1385),
    .A1(\vmem[292] ),
    .S(_06726_),
    .X(_01859_));
 or4_1 _22471_ (.A(net721),
    .B(net641),
    .C(net853),
    .D(_06496_),
    .X(_06727_));
 mux2_1 _22472_ (.A0(net1330),
    .A1(\vmem[291] ),
    .S(_06727_),
    .X(_01860_));
 or4_1 _22473_ (.A(net744),
    .B(net663),
    .C(net875),
    .D(_06499_),
    .X(_06728_));
 mux2_1 _22474_ (.A0(net1373),
    .A1(\vmem[290] ),
    .S(_06728_),
    .X(_01861_));
 or4_1 _22475_ (.A(net746),
    .B(net666),
    .C(net877),
    .D(_06502_),
    .X(_06729_));
 mux2_1 _22476_ (.A0(net1376),
    .A1(\vmem[289] ),
    .S(_06729_),
    .X(_01862_));
 or4_1 _22477_ (.A(net728),
    .B(net646),
    .C(net860),
    .D(_06505_),
    .X(_06730_));
 mux2_1 _22478_ (.A0(net1342),
    .A1(\vmem[288] ),
    .S(_06730_),
    .X(_01863_));
 or4_1 _22479_ (.A(net735),
    .B(net655),
    .C(net866),
    .D(_06507_),
    .X(_06731_));
 mux2_1 _22480_ (.A0(net1356),
    .A1(\vmem[287] ),
    .S(_06731_),
    .X(_01864_));
 or4_1 _22481_ (.A(net740),
    .B(net660),
    .C(net870),
    .D(_06509_),
    .X(_06732_));
 mux2_1 _22482_ (.A0(net1369),
    .A1(\vmem[286] ),
    .S(_06732_),
    .X(_01865_));
 or4_1 _22483_ (.A(net739),
    .B(net661),
    .C(net872),
    .D(_06511_),
    .X(_06733_));
 mux2_1 _22484_ (.A0(net1364),
    .A1(\vmem[285] ),
    .S(_06733_),
    .X(_01866_));
 or4_1 _22485_ (.A(net756),
    .B(net671),
    .C(net881),
    .D(_06513_),
    .X(_06734_));
 mux2_1 _22486_ (.A0(net1388),
    .A1(\vmem[284] ),
    .S(_06734_),
    .X(_01867_));
 or4_1 _22487_ (.A(net737),
    .B(net657),
    .C(net868),
    .D(_06515_),
    .X(_06735_));
 mux2_1 _22488_ (.A0(net1362),
    .A1(\vmem[283] ),
    .S(_06735_),
    .X(_01868_));
 or4_1 _22489_ (.A(net731),
    .B(net650),
    .C(net863),
    .D(_06517_),
    .X(_06736_));
 mux2_1 _22490_ (.A0(net1347),
    .A1(\vmem[282] ),
    .S(_06736_),
    .X(_01869_));
 or4_1 _22491_ (.A(net733),
    .B(net652),
    .C(net865),
    .D(_06519_),
    .X(_06737_));
 mux2_1 _22492_ (.A0(net1351),
    .A1(\vmem[281] ),
    .S(_06737_),
    .X(_01870_));
 or4_1 _22493_ (.A(net725),
    .B(net643),
    .C(net857),
    .D(_06521_),
    .X(_06738_));
 mux2_1 _22494_ (.A0(net1338),
    .A1(\vmem[280] ),
    .S(_06738_),
    .X(_01871_));
 or4_1 _22495_ (.A(net732),
    .B(net651),
    .C(net862),
    .D(_06523_),
    .X(_06739_));
 mux2_1 _22496_ (.A0(net1349),
    .A1(\vmem[279] ),
    .S(_06739_),
    .X(_01872_));
 or4_1 _22497_ (.A(net754),
    .B(net674),
    .C(net883),
    .D(_06525_),
    .X(_06740_));
 mux2_1 _22498_ (.A0(net1390),
    .A1(\vmem[278] ),
    .S(_06740_),
    .X(_01873_));
 or4_1 _22499_ (.A(net727),
    .B(net645),
    .C(net856),
    .D(_06527_),
    .X(_06741_));
 mux2_1 _22500_ (.A0(net1340),
    .A1(\vmem[277] ),
    .S(_06741_),
    .X(_01874_));
 or4_1 _22501_ (.A(net751),
    .B(net669),
    .C(net885),
    .D(_06529_),
    .X(_06742_));
 mux2_1 _22502_ (.A0(net1384),
    .A1(\vmem[276] ),
    .S(_06742_),
    .X(_01875_));
 or4_1 _22503_ (.A(net721),
    .B(net641),
    .C(net854),
    .D(_06531_),
    .X(_06743_));
 mux2_1 _22504_ (.A0(net1330),
    .A1(\vmem[275] ),
    .S(_06743_),
    .X(_01876_));
 or4_1 _22505_ (.A(net744),
    .B(net663),
    .C(net875),
    .D(_06533_),
    .X(_06744_));
 mux2_1 _22506_ (.A0(net1373),
    .A1(\vmem[274] ),
    .S(_06744_),
    .X(_01877_));
 or4_1 _22507_ (.A(net746),
    .B(net666),
    .C(net877),
    .D(_06535_),
    .X(_06745_));
 mux2_1 _22508_ (.A0(net1376),
    .A1(\vmem[273] ),
    .S(_06745_),
    .X(_01878_));
 or4_1 _22509_ (.A(net727),
    .B(net645),
    .C(net859),
    .D(_06537_),
    .X(_06746_));
 mux2_1 _22510_ (.A0(net1340),
    .A1(\vmem[272] ),
    .S(_06746_),
    .X(_01879_));
 or4_1 _22511_ (.A(net735),
    .B(net655),
    .C(net866),
    .D(_06539_),
    .X(_06747_));
 mux2_1 _22512_ (.A0(net1356),
    .A1(\vmem[271] ),
    .S(_06747_),
    .X(_01880_));
 or4_1 _22513_ (.A(net740),
    .B(net660),
    .C(net870),
    .D(_06541_),
    .X(_06748_));
 mux2_1 _22514_ (.A0(net1367),
    .A1(\vmem[270] ),
    .S(_06748_),
    .X(_01881_));
 or4_1 _22515_ (.A(net736),
    .B(net656),
    .C(net867),
    .D(_06543_),
    .X(_06749_));
 mux2_1 _22516_ (.A0(net1359),
    .A1(\vmem[269] ),
    .S(_06749_),
    .X(_01882_));
 or4_1 _22517_ (.A(net756),
    .B(net671),
    .C(net882),
    .D(_06545_),
    .X(_06750_));
 mux2_1 _22518_ (.A0(net1388),
    .A1(\vmem[268] ),
    .S(_06750_),
    .X(_01883_));
 or4_1 _22519_ (.A(net737),
    .B(net657),
    .C(net868),
    .D(_06547_),
    .X(_06751_));
 mux2_1 _22520_ (.A0(net1360),
    .A1(\vmem[267] ),
    .S(_06751_),
    .X(_01884_));
 or4_1 _22521_ (.A(net731),
    .B(net650),
    .C(net863),
    .D(_06549_),
    .X(_06752_));
 mux2_1 _22522_ (.A0(net1347),
    .A1(\vmem[266] ),
    .S(_06752_),
    .X(_01885_));
 or4_1 _22523_ (.A(net744),
    .B(net663),
    .C(net874),
    .D(_06551_),
    .X(_06753_));
 mux2_1 _22524_ (.A0(net1373),
    .A1(\vmem[265] ),
    .S(_06753_),
    .X(_01886_));
 or4_1 _22525_ (.A(net726),
    .B(net644),
    .C(net858),
    .D(_06553_),
    .X(_06754_));
 mux2_1 _22526_ (.A0(net1343),
    .A1(\vmem[264] ),
    .S(_06754_),
    .X(_01887_));
 or4_1 _22527_ (.A(net734),
    .B(net652),
    .C(net865),
    .D(_06555_),
    .X(_06755_));
 mux2_1 _22528_ (.A0(net1352),
    .A1(\vmem[263] ),
    .S(_06755_),
    .X(_01888_));
 or4_1 _22529_ (.A(net754),
    .B(net672),
    .C(net881),
    .D(_06557_),
    .X(_06756_));
 mux2_1 _22530_ (.A0(net1391),
    .A1(\vmem[262] ),
    .S(_06756_),
    .X(_01889_));
 or4_1 _22531_ (.A(net724),
    .B(net644),
    .C(net855),
    .D(_06559_),
    .X(_06757_));
 mux2_1 _22532_ (.A0(net1336),
    .A1(\vmem[261] ),
    .S(_06757_),
    .X(_01890_));
 or4_1 _22533_ (.A(net751),
    .B(net669),
    .C(net879),
    .D(_06561_),
    .X(_06758_));
 mux2_1 _22534_ (.A0(net1384),
    .A1(\vmem[260] ),
    .S(_06758_),
    .X(_01891_));
 or4_1 _22535_ (.A(net721),
    .B(net641),
    .C(net854),
    .D(_06563_),
    .X(_06759_));
 mux2_1 _22536_ (.A0(net1332),
    .A1(\vmem[259] ),
    .S(_06759_),
    .X(_01892_));
 or4_1 _22537_ (.A(net744),
    .B(net663),
    .C(net875),
    .D(_06565_),
    .X(_06760_));
 mux2_1 _22538_ (.A0(net1373),
    .A1(\vmem[258] ),
    .S(_06760_),
    .X(_01893_));
 or4_1 _22539_ (.A(net746),
    .B(net666),
    .C(net877),
    .D(_06567_),
    .X(_06761_));
 mux2_1 _22540_ (.A0(net1376),
    .A1(\vmem[257] ),
    .S(_06761_),
    .X(_01894_));
 or4_1 _22541_ (.A(net727),
    .B(net645),
    .C(net859),
    .D(_06569_),
    .X(_06762_));
 mux2_1 _22542_ (.A0(net1340),
    .A1(\vmem[256] ),
    .S(_06762_),
    .X(_01895_));
 o21ai_4 _22543_ (.A1(\stadly_mpw03_prog_rise_9.Y ),
    .A2(net1327),
    .B1(_09415_),
    .Y(_06763_));
 or4_1 _22544_ (.A(net773),
    .B(net615),
    .C(_06410_),
    .D(net832),
    .X(_06764_));
 mux2_1 _22545_ (.A0(net1349),
    .A1(\vmem[255] ),
    .S(_06764_),
    .X(_01896_));
 or4_1 _22546_ (.A(net783),
    .B(net622),
    .C(_06414_),
    .D(net839),
    .X(_06765_));
 mux2_1 _22547_ (.A0(net1368),
    .A1(\vmem[254] ),
    .S(_06765_),
    .X(_01897_));
 or4_1 _22548_ (.A(net781),
    .B(net623),
    .C(_06417_),
    .D(net838),
    .X(_06766_));
 mux2_1 _22549_ (.A0(net1365),
    .A1(\vmem[253] ),
    .S(_06766_),
    .X(_01898_));
 or4_1 _22550_ (.A(net789),
    .B(net627),
    .C(_06420_),
    .D(net844),
    .X(_06767_));
 mux2_1 _22551_ (.A0(net1376),
    .A1(\vmem[252] ),
    .S(_06767_),
    .X(_01899_));
 or4_1 _22552_ (.A(net779),
    .B(net624),
    .C(_06423_),
    .D(net835),
    .X(_06768_));
 mux2_1 _22553_ (.A0(net1360),
    .A1(\vmem[251] ),
    .S(_06768_),
    .X(_01900_));
 or4_1 _22554_ (.A(net765),
    .B(net611),
    .C(_06426_),
    .D(net826),
    .X(_06769_));
 mux2_1 _22555_ (.A0(net1339),
    .A1(\vmem[250] ),
    .S(_06769_),
    .X(_01901_));
 or4_1 _22556_ (.A(net786),
    .B(net625),
    .C(_06429_),
    .D(net842),
    .X(_06770_));
 mux2_1 _22557_ (.A0(net1351),
    .A1(\vmem[249] ),
    .S(_06770_),
    .X(_01902_));
 or4_1 _22558_ (.A(net763),
    .B(net609),
    .C(_06432_),
    .D(net824),
    .X(_06771_));
 mux2_1 _22559_ (.A0(net1335),
    .A1(\vmem[248] ),
    .S(_06771_),
    .X(_01903_));
 or4_1 _22560_ (.A(net775),
    .B(net617),
    .C(_06435_),
    .D(net834),
    .X(_06772_));
 mux2_1 _22561_ (.A0(net1353),
    .A1(\vmem[247] ),
    .S(_06772_),
    .X(_01904_));
 or4_1 _22562_ (.A(net793),
    .B(net636),
    .C(_06438_),
    .D(net848),
    .X(_06773_));
 mux2_1 _22563_ (.A0(net1384),
    .A1(\vmem[246] ),
    .S(_06773_),
    .X(_01905_));
 or4_1 _22564_ (.A(net761),
    .B(net605),
    .C(_06441_),
    .D(net822),
    .X(_06774_));
 mux2_1 _22565_ (.A0(net1331),
    .A1(\vmem[245] ),
    .S(_06774_),
    .X(_01906_));
 or4_1 _22566_ (.A(net793),
    .B(net631),
    .C(_06444_),
    .D(net847),
    .X(_06775_));
 mux2_1 _22567_ (.A0(net1383),
    .A1(\vmem[244] ),
    .S(_06775_),
    .X(_01907_));
 or4_1 _22568_ (.A(net758),
    .B(net604),
    .C(_06447_),
    .D(net820),
    .X(_06776_));
 mux2_1 _22569_ (.A0(net1327),
    .A1(\vmem[243] ),
    .S(_06776_),
    .X(_01908_));
 or4_1 _22570_ (.A(net787),
    .B(net626),
    .C(_06450_),
    .D(net843),
    .X(_06777_));
 mux2_1 _22571_ (.A0(net1374),
    .A1(\vmem[242] ),
    .S(_06777_),
    .X(_01909_));
 or4_1 _22572_ (.A(net791),
    .B(net629),
    .C(_06453_),
    .D(net845),
    .X(_06778_));
 mux2_1 _22573_ (.A0(net1379),
    .A1(\vmem[241] ),
    .S(_06778_),
    .X(_01910_));
 or4_1 _22574_ (.A(net762),
    .B(net606),
    .C(_06457_),
    .D(net823),
    .X(_06779_));
 mux2_1 _22575_ (.A0(net1333),
    .A1(\vmem[240] ),
    .S(_06779_),
    .X(_01911_));
 or4_1 _22576_ (.A(net772),
    .B(net615),
    .C(_06460_),
    .D(net832),
    .X(_06780_));
 mux2_1 _22577_ (.A0(net1348),
    .A1(\vmem[239] ),
    .S(_06780_),
    .X(_01912_));
 or4_1 _22578_ (.A(net783),
    .B(net622),
    .C(_06463_),
    .D(net840),
    .X(_06781_));
 mux2_1 _22579_ (.A0(net1368),
    .A1(\vmem[238] ),
    .S(_06781_),
    .X(_01913_));
 or4_1 _22580_ (.A(net784),
    .B(net630),
    .C(_06466_),
    .D(net840),
    .X(_06782_));
 mux2_1 _22581_ (.A0(net1382),
    .A1(\vmem[237] ),
    .S(_06782_),
    .X(_01914_));
 or4_1 _22582_ (.A(net789),
    .B(net627),
    .C(_06469_),
    .D(net844),
    .X(_06783_));
 mux2_1 _22583_ (.A0(net1378),
    .A1(\vmem[236] ),
    .S(_06783_),
    .X(_01915_));
 or4_1 _22584_ (.A(net779),
    .B(net620),
    .C(_06472_),
    .D(net835),
    .X(_06784_));
 mux2_1 _22585_ (.A0(net1361),
    .A1(\vmem[235] ),
    .S(_06784_),
    .X(_01916_));
 or4_1 _22586_ (.A(net765),
    .B(net611),
    .C(_06475_),
    .D(net826),
    .X(_06785_));
 mux2_1 _22587_ (.A0(net1339),
    .A1(\vmem[234] ),
    .S(_06785_),
    .X(_01917_));
 or4_1 _22588_ (.A(net786),
    .B(net625),
    .C(_06478_),
    .D(net842),
    .X(_06786_));
 mux2_1 _22589_ (.A0(net1371),
    .A1(\vmem[233] ),
    .S(_06786_),
    .X(_01918_));
 or4_1 _22590_ (.A(net763),
    .B(net609),
    .C(_06481_),
    .D(net824),
    .X(_06787_));
 mux2_1 _22591_ (.A0(net1337),
    .A1(\vmem[232] ),
    .S(_06787_),
    .X(_01919_));
 or4_1 _22592_ (.A(net775),
    .B(net617),
    .C(_06484_),
    .D(net834),
    .X(_06788_));
 mux2_1 _22593_ (.A0(net1353),
    .A1(\vmem[231] ),
    .S(_06788_),
    .X(_01920_));
 or4_1 _22594_ (.A(net797),
    .B(net636),
    .C(_06487_),
    .D(net849),
    .X(_06789_));
 mux2_1 _22595_ (.A0(net1390),
    .A1(\vmem[230] ),
    .S(_06789_),
    .X(_01921_));
 or4_1 _22596_ (.A(net761),
    .B(net605),
    .C(_06490_),
    .D(net822),
    .X(_06790_));
 mux2_1 _22597_ (.A0(net1331),
    .A1(\vmem[229] ),
    .S(_06790_),
    .X(_01922_));
 or4_1 _22598_ (.A(net793),
    .B(net631),
    .C(_06493_),
    .D(net848),
    .X(_06791_));
 mux2_1 _22599_ (.A0(net1385),
    .A1(\vmem[228] ),
    .S(_06791_),
    .X(_01923_));
 or4_1 _22600_ (.A(net758),
    .B(net604),
    .C(_06496_),
    .D(net820),
    .X(_06792_));
 mux2_1 _22601_ (.A0(net1328),
    .A1(\vmem[227] ),
    .S(_06792_),
    .X(_01924_));
 or4_1 _22602_ (.A(net787),
    .B(net626),
    .C(_06499_),
    .D(net843),
    .X(_06793_));
 mux2_1 _22603_ (.A0(net1374),
    .A1(\vmem[226] ),
    .S(_06793_),
    .X(_01925_));
 or4_1 _22604_ (.A(net791),
    .B(net629),
    .C(_06502_),
    .D(net844),
    .X(_06794_));
 mux2_1 _22605_ (.A0(net1379),
    .A1(\vmem[225] ),
    .S(_06794_),
    .X(_01926_));
 or4_1 _22606_ (.A(net762),
    .B(net606),
    .C(_06505_),
    .D(net823),
    .X(_06795_));
 mux2_1 _22607_ (.A0(net1333),
    .A1(\vmem[224] ),
    .S(_06795_),
    .X(_01927_));
 or4_1 _22608_ (.A(net773),
    .B(net615),
    .C(_06507_),
    .D(net832),
    .X(_06796_));
 mux2_1 _22609_ (.A0(net1349),
    .A1(\vmem[223] ),
    .S(_06796_),
    .X(_01928_));
 or4_1 _22610_ (.A(net782),
    .B(net623),
    .C(_06509_),
    .D(net839),
    .X(_06797_));
 mux2_1 _22611_ (.A0(net1364),
    .A1(\vmem[222] ),
    .S(_06797_),
    .X(_01929_));
 or4_1 _22612_ (.A(net784),
    .B(net621),
    .C(_06511_),
    .D(net838),
    .X(_06798_));
 mux2_1 _22613_ (.A0(net1365),
    .A1(\vmem[221] ),
    .S(_06798_),
    .X(_01930_));
 or4_1 _22614_ (.A(net795),
    .B(net634),
    .C(_06513_),
    .D(net846),
    .X(_06799_));
 mux2_1 _22615_ (.A0(net1381),
    .A1(\vmem[220] ),
    .S(_06799_),
    .X(_01931_));
 or4_1 _22616_ (.A(net778),
    .B(net619),
    .C(_06515_),
    .D(net836),
    .X(_06800_));
 mux2_1 _22617_ (.A0(net1359),
    .A1(\vmem[219] ),
    .S(_06800_),
    .X(_01932_));
 or4_1 _22618_ (.A(net770),
    .B(net614),
    .C(_06517_),
    .D(net830),
    .X(_06801_));
 mux2_1 _22619_ (.A0(net1345),
    .A1(\vmem[218] ),
    .S(_06801_),
    .X(_01933_));
 or4_1 _22620_ (.A(net767),
    .B(net612),
    .C(_06519_),
    .D(net833),
    .X(_06802_));
 mux2_1 _22621_ (.A0(net1355),
    .A1(\vmem[217] ),
    .S(_06802_),
    .X(_01934_));
 or4_1 _22622_ (.A(net763),
    .B(net609),
    .C(_06521_),
    .D(net824),
    .X(_06803_));
 mux2_1 _22623_ (.A0(net1335),
    .A1(\vmem[216] ),
    .S(_06803_),
    .X(_01935_));
 or4_1 _22624_ (.A(net774),
    .B(net616),
    .C(_06523_),
    .D(net834),
    .X(_06804_));
 mux2_1 _22625_ (.A0(net1352),
    .A1(\vmem[215] ),
    .S(_06804_),
    .X(_01936_));
 or4_1 _22626_ (.A(net796),
    .B(net635),
    .C(_06525_),
    .D(net850),
    .X(_06805_));
 mux2_1 _22627_ (.A0(net1389),
    .A1(\vmem[214] ),
    .S(_06805_),
    .X(_01937_));
 or4_1 _22628_ (.A(net763),
    .B(net609),
    .C(_06527_),
    .D(net824),
    .X(_06806_));
 mux2_1 _22629_ (.A0(net1335),
    .A1(\vmem[213] ),
    .S(_06806_),
    .X(_01938_));
 or4_1 _22630_ (.A(net793),
    .B(net631),
    .C(_06529_),
    .D(net847),
    .X(_06807_));
 mux2_1 _22631_ (.A0(net1383),
    .A1(\vmem[212] ),
    .S(_06807_),
    .X(_01939_));
 or4_1 _22632_ (.A(net758),
    .B(net604),
    .C(_06531_),
    .D(net820),
    .X(_06808_));
 mux2_1 _22633_ (.A0(net1327),
    .A1(\vmem[211] ),
    .S(_06808_),
    .X(_01940_));
 or4_1 _22634_ (.A(net787),
    .B(net626),
    .C(_06533_),
    .D(net843),
    .X(_06809_));
 mux2_1 _22635_ (.A0(net1374),
    .A1(\vmem[210] ),
    .S(_06809_),
    .X(_01941_));
 or4_1 _22636_ (.A(net789),
    .B(net627),
    .C(_06535_),
    .D(net844),
    .X(_06810_));
 mux2_1 _22637_ (.A0(net1376),
    .A1(\vmem[209] ),
    .S(_06810_),
    .X(_01942_));
 or4_1 _22638_ (.A(net766),
    .B(net612),
    .C(_06537_),
    .D(net827),
    .X(_06811_));
 mux2_1 _22639_ (.A0(net1340),
    .A1(\vmem[208] ),
    .S(_06811_),
    .X(_01943_));
 or4_1 _22640_ (.A(net778),
    .B(net618),
    .C(_06539_),
    .D(net836),
    .X(_06812_));
 mux2_1 _22641_ (.A0(net1358),
    .A1(\vmem[207] ),
    .S(_06812_),
    .X(_01944_));
 or4_1 _22642_ (.A(net781),
    .B(net621),
    .C(_06541_),
    .D(net838),
    .X(_06813_));
 mux2_1 _22643_ (.A0(net1366),
    .A1(\vmem[206] ),
    .S(_06813_),
    .X(_01945_));
 or4_1 _22644_ (.A(net784),
    .B(net621),
    .C(_06543_),
    .D(net838),
    .X(_06814_));
 mux2_1 _22645_ (.A0(net1366),
    .A1(\vmem[205] ),
    .S(_06814_),
    .X(_01946_));
 or4_1 _22646_ (.A(net796),
    .B(net634),
    .C(_06545_),
    .D(net850),
    .X(_06815_));
 mux2_1 _22647_ (.A0(net1386),
    .A1(\vmem[204] ),
    .S(_06815_),
    .X(_01947_));
 or4_1 _22648_ (.A(net777),
    .B(net618),
    .C(_06547_),
    .D(net837),
    .X(_06816_));
 mux2_1 _22649_ (.A0(net1358),
    .A1(\vmem[203] ),
    .S(_06816_),
    .X(_01948_));
 or4_1 _22650_ (.A(net770),
    .B(net614),
    .C(_06549_),
    .D(net830),
    .X(_06817_));
 mux2_1 _22651_ (.A0(net1345),
    .A1(\vmem[202] ),
    .S(_06817_),
    .X(_01949_));
 or4_1 _22652_ (.A(net767),
    .B(net613),
    .C(_06551_),
    .D(net828),
    .X(_06818_));
 mux2_1 _22653_ (.A0(net1355),
    .A1(\vmem[201] ),
    .S(_06818_),
    .X(_01950_));
 or4_1 _22654_ (.A(net763),
    .B(net609),
    .C(_06553_),
    .D(net824),
    .X(_06819_));
 mux2_1 _22655_ (.A0(net1335),
    .A1(\vmem[200] ),
    .S(_06819_),
    .X(_01951_));
 or4_1 _22656_ (.A(net775),
    .B(net616),
    .C(_06555_),
    .D(net833),
    .X(_06820_));
 mux2_1 _22657_ (.A0(net1353),
    .A1(\vmem[199] ),
    .S(_06820_),
    .X(_01952_));
 or4_1 _22658_ (.A(net796),
    .B(net634),
    .C(_06557_),
    .D(net849),
    .X(_06821_));
 mux2_1 _22659_ (.A0(net1389),
    .A1(\vmem[198] ),
    .S(_06821_),
    .X(_01953_));
 or4_1 _22660_ (.A(net764),
    .B(net610),
    .C(_06559_),
    .D(net825),
    .X(_06822_));
 mux2_1 _22661_ (.A0(net1336),
    .A1(\vmem[197] ),
    .S(_06822_),
    .X(_01954_));
 or4_1 _22662_ (.A(net793),
    .B(net631),
    .C(_06561_),
    .D(net847),
    .X(_06823_));
 mux2_1 _22663_ (.A0(net1383),
    .A1(\vmem[196] ),
    .S(_06823_),
    .X(_01955_));
 or4_1 _22664_ (.A(net758),
    .B(net604),
    .C(_06563_),
    .D(net820),
    .X(_06824_));
 mux2_1 _22665_ (.A0(net1327),
    .A1(\vmem[195] ),
    .S(_06824_),
    .X(_01956_));
 or4_1 _22666_ (.A(net787),
    .B(net626),
    .C(_06565_),
    .D(net843),
    .X(_06825_));
 mux2_1 _22667_ (.A0(net1374),
    .A1(\vmem[194] ),
    .S(_06825_),
    .X(_01957_));
 or4_1 _22668_ (.A(net789),
    .B(net627),
    .C(_06567_),
    .D(net844),
    .X(_06826_));
 mux2_1 _22669_ (.A0(net1376),
    .A1(\vmem[193] ),
    .S(_06826_),
    .X(_01958_));
 or4_1 _22670_ (.A(net762),
    .B(net606),
    .C(_06569_),
    .D(net823),
    .X(_06827_));
 mux2_1 _22671_ (.A0(net1333),
    .A1(\vmem[192] ),
    .S(_06827_),
    .X(_01959_));
 or4_1 _22672_ (.A(net735),
    .B(net619),
    .C(_06410_),
    .D(net836),
    .X(_06828_));
 mux2_1 _22673_ (.A0(net1356),
    .A1(\vmem[191] ),
    .S(_06828_),
    .X(_01960_));
 or4_1 _22674_ (.A(net741),
    .B(net622),
    .C(_06414_),
    .D(net839),
    .X(_06829_));
 mux2_1 _22675_ (.A0(net1366),
    .A1(\vmem[190] ),
    .S(_06829_),
    .X(_01961_));
 or4_1 _22676_ (.A(net739),
    .B(net621),
    .C(_06417_),
    .D(net838),
    .X(_06830_));
 mux2_1 _22677_ (.A0(net1365),
    .A1(\vmem[189] ),
    .S(_06830_),
    .X(_01962_));
 or4_1 _22678_ (.A(net746),
    .B(net627),
    .C(_06420_),
    .D(net844),
    .X(_06831_));
 mux2_1 _22679_ (.A0(net1376),
    .A1(\vmem[188] ),
    .S(_06831_),
    .X(_01963_));
 or4_1 _22680_ (.A(net737),
    .B(net620),
    .C(_06423_),
    .D(net837),
    .X(_06832_));
 mux2_1 _22681_ (.A0(net1361),
    .A1(\vmem[187] ),
    .S(_06832_),
    .X(_01964_));
 or4_1 _22682_ (.A(net725),
    .B(net611),
    .C(_06426_),
    .D(net826),
    .X(_06833_));
 mux2_1 _22683_ (.A0(net1338),
    .A1(\vmem[186] ),
    .S(_06833_),
    .X(_01965_));
 or4_1 _22684_ (.A(net743),
    .B(net625),
    .C(_06429_),
    .D(net842),
    .X(_06834_));
 mux2_1 _22685_ (.A0(net1371),
    .A1(\vmem[185] ),
    .S(_06834_),
    .X(_01966_));
 or4_1 _22686_ (.A(net724),
    .B(net609),
    .C(_06432_),
    .D(net824),
    .X(_06835_));
 mux2_1 _22687_ (.A0(net1335),
    .A1(\vmem[184] ),
    .S(_06835_),
    .X(_01967_));
 or4_1 _22688_ (.A(net733),
    .B(net617),
    .C(_06435_),
    .D(net833),
    .X(_06836_));
 mux2_1 _22689_ (.A0(net1355),
    .A1(\vmem[183] ),
    .S(_06836_),
    .X(_01968_));
 or4_1 _22690_ (.A(net755),
    .B(net636),
    .C(_06438_),
    .D(net849),
    .X(_06837_));
 mux2_1 _22691_ (.A0(net1390),
    .A1(\vmem[182] ),
    .S(_06837_),
    .X(_01969_));
 or4_1 _22692_ (.A(net722),
    .B(net608),
    .C(_06441_),
    .D(net822),
    .X(_06838_));
 mux2_1 _22693_ (.A0(net1332),
    .A1(\vmem[181] ),
    .S(_06838_),
    .X(_01970_));
 or4_1 _22694_ (.A(net750),
    .B(net632),
    .C(_06444_),
    .D(net847),
    .X(_06839_));
 mux2_1 _22695_ (.A0(net1385),
    .A1(\vmem[180] ),
    .S(_06839_),
    .X(_01971_));
 or4_1 _22696_ (.A(net720),
    .B(net604),
    .C(_06447_),
    .D(net820),
    .X(_06840_));
 mux2_1 _22697_ (.A0(net1327),
    .A1(\vmem[179] ),
    .S(_06840_),
    .X(_01972_));
 or4_1 _22698_ (.A(net744),
    .B(net626),
    .C(_06450_),
    .D(net843),
    .X(_06841_));
 mux2_1 _22699_ (.A0(net1373),
    .A1(\vmem[178] ),
    .S(_06841_),
    .X(_01973_));
 or4_1 _22700_ (.A(net748),
    .B(net629),
    .C(_06453_),
    .D(net845),
    .X(_06842_));
 mux2_1 _22701_ (.A0(net1379),
    .A1(\vmem[177] ),
    .S(_06842_),
    .X(_01974_));
 or4_1 _22702_ (.A(net723),
    .B(net607),
    .C(_06457_),
    .D(net823),
    .X(_06843_));
 mux2_1 _22703_ (.A0(net1334),
    .A1(\vmem[176] ),
    .S(_06843_),
    .X(_01975_));
 or4_1 _22704_ (.A(net731),
    .B(net615),
    .C(_06460_),
    .D(net832),
    .X(_06844_));
 mux2_1 _22705_ (.A0(net1348),
    .A1(\vmem[175] ),
    .S(_06844_),
    .X(_01976_));
 or4_1 _22706_ (.A(net750),
    .B(net631),
    .C(_06463_),
    .D(net847),
    .X(_06845_));
 mux2_1 _22707_ (.A0(net1368),
    .A1(\vmem[174] ),
    .S(_06845_),
    .X(_01977_));
 or4_1 _22708_ (.A(net742),
    .B(net621),
    .C(_06466_),
    .D(net840),
    .X(_06846_));
 mux2_1 _22709_ (.A0(net1365),
    .A1(\vmem[173] ),
    .S(_06846_),
    .X(_01978_));
 or4_1 _22710_ (.A(net746),
    .B(net627),
    .C(_06469_),
    .D(net844),
    .X(_06847_));
 mux2_1 _22711_ (.A0(net1376),
    .A1(\vmem[172] ),
    .S(_06847_),
    .X(_01979_));
 or4_1 _22712_ (.A(net738),
    .B(net620),
    .C(_06472_),
    .D(net837),
    .X(_06848_));
 mux2_1 _22713_ (.A0(net1361),
    .A1(\vmem[171] ),
    .S(_06848_),
    .X(_01980_));
 or4_1 _22714_ (.A(net725),
    .B(net611),
    .C(_06475_),
    .D(net828),
    .X(_06849_));
 mux2_1 _22715_ (.A0(net1339),
    .A1(\vmem[170] ),
    .S(_06849_),
    .X(_01981_));
 or4_1 _22716_ (.A(net743),
    .B(net625),
    .C(_06478_),
    .D(net842),
    .X(_06850_));
 mux2_1 _22717_ (.A0(net1371),
    .A1(\vmem[169] ),
    .S(_06850_),
    .X(_01982_));
 or4_1 _22718_ (.A(net724),
    .B(net609),
    .C(_06481_),
    .D(net824),
    .X(_06851_));
 mux2_1 _22719_ (.A0(net1335),
    .A1(\vmem[168] ),
    .S(_06851_),
    .X(_01983_));
 or4_1 _22720_ (.A(net733),
    .B(net617),
    .C(_06484_),
    .D(net833),
    .X(_06852_));
 mux2_1 _22721_ (.A0(net1351),
    .A1(\vmem[167] ),
    .S(_06852_),
    .X(_01984_));
 or4_1 _22722_ (.A(net755),
    .B(net636),
    .C(_06487_),
    .D(net849),
    .X(_06853_));
 mux2_1 _22723_ (.A0(net1390),
    .A1(\vmem[166] ),
    .S(_06853_),
    .X(_01985_));
 or4_1 _22724_ (.A(net722),
    .B(net605),
    .C(_06490_),
    .D(net822),
    .X(_06854_));
 mux2_1 _22725_ (.A0(net1331),
    .A1(\vmem[165] ),
    .S(_06854_),
    .X(_01986_));
 or4_1 _22726_ (.A(net750),
    .B(net631),
    .C(_06493_),
    .D(net847),
    .X(_06855_));
 mux2_1 _22727_ (.A0(net1383),
    .A1(\vmem[164] ),
    .S(_06855_),
    .X(_01987_));
 or4_1 _22728_ (.A(net720),
    .B(net604),
    .C(_06496_),
    .D(net821),
    .X(_06856_));
 mux2_1 _22729_ (.A0(net1328),
    .A1(\vmem[163] ),
    .S(_06856_),
    .X(_01988_));
 or4_1 _22730_ (.A(net744),
    .B(net626),
    .C(_06499_),
    .D(net843),
    .X(_06857_));
 mux2_1 _22731_ (.A0(net1373),
    .A1(\vmem[162] ),
    .S(_06857_),
    .X(_01989_));
 or4_1 _22732_ (.A(net748),
    .B(net629),
    .C(_06502_),
    .D(net845),
    .X(_06858_));
 mux2_1 _22733_ (.A0(net1379),
    .A1(\vmem[161] ),
    .S(_06858_),
    .X(_01990_));
 or4_1 _22734_ (.A(net723),
    .B(net606),
    .C(_06505_),
    .D(net823),
    .X(_06859_));
 mux2_1 _22735_ (.A0(net1334),
    .A1(\vmem[160] ),
    .S(_06859_),
    .X(_01991_));
 or4_1 _22736_ (.A(net731),
    .B(net615),
    .C(_06507_),
    .D(net832),
    .X(_06860_));
 mux2_1 _22737_ (.A0(net1349),
    .A1(\vmem[159] ),
    .S(_06860_),
    .X(_01992_));
 or4_1 _22738_ (.A(net741),
    .B(net622),
    .C(_06509_),
    .D(net840),
    .X(_06861_));
 mux2_1 _22739_ (.A0(net1368),
    .A1(\vmem[158] ),
    .S(_06861_),
    .X(_01993_));
 or4_1 _22740_ (.A(net739),
    .B(net621),
    .C(_06511_),
    .D(net838),
    .X(_06862_));
 mux2_1 _22741_ (.A0(net1365),
    .A1(\vmem[157] ),
    .S(_06862_),
    .X(_01994_));
 or4_1 _22742_ (.A(net753),
    .B(net634),
    .C(_06513_),
    .D(net846),
    .X(_06863_));
 mux2_1 _22743_ (.A0(net1381),
    .A1(\vmem[156] ),
    .S(_06863_),
    .X(_01995_));
 or4_1 _22744_ (.A(net735),
    .B(net618),
    .C(_06515_),
    .D(net836),
    .X(_06864_));
 mux2_1 _22745_ (.A0(net1359),
    .A1(\vmem[155] ),
    .S(_06864_),
    .X(_01996_));
 or4_1 _22746_ (.A(net730),
    .B(net614),
    .C(_06517_),
    .D(net830),
    .X(_06865_));
 mux2_1 _22747_ (.A0(net1345),
    .A1(\vmem[154] ),
    .S(_06865_),
    .X(_01997_));
 or4_1 _22748_ (.A(net727),
    .B(net613),
    .C(_06519_),
    .D(net827),
    .X(_06866_));
 mux2_1 _22749_ (.A0(net1342),
    .A1(\vmem[153] ),
    .S(_06866_),
    .X(_01998_));
 or4_1 _22750_ (.A(net724),
    .B(net609),
    .C(_06521_),
    .D(net824),
    .X(_06867_));
 mux2_1 _22751_ (.A0(net1335),
    .A1(\vmem[152] ),
    .S(_06867_),
    .X(_01999_));
 or4_1 _22752_ (.A(net733),
    .B(net617),
    .C(_06523_),
    .D(net833),
    .X(_06868_));
 mux2_1 _22753_ (.A0(net1351),
    .A1(\vmem[151] ),
    .S(_06868_),
    .X(_02000_));
 or4_1 _22754_ (.A(net753),
    .B(net634),
    .C(_06525_),
    .D(net849),
    .X(_06869_));
 mux2_1 _22755_ (.A0(net1386),
    .A1(\vmem[150] ),
    .S(_06869_),
    .X(_02001_));
 or4_1 _22756_ (.A(net721),
    .B(net605),
    .C(_06527_),
    .D(net823),
    .X(_06870_));
 mux2_1 _22757_ (.A0(net1332),
    .A1(\vmem[149] ),
    .S(_06870_),
    .X(_02002_));
 or4_1 _22758_ (.A(net750),
    .B(net631),
    .C(_06529_),
    .D(net847),
    .X(_06871_));
 mux2_1 _22759_ (.A0(net1385),
    .A1(\vmem[148] ),
    .S(_06871_),
    .X(_02003_));
 or4_1 _22760_ (.A(net720),
    .B(net604),
    .C(_06531_),
    .D(net820),
    .X(_06872_));
 mux2_1 _22761_ (.A0(net1327),
    .A1(\vmem[147] ),
    .S(_06872_),
    .X(_02004_));
 or4_1 _22762_ (.A(net744),
    .B(net626),
    .C(_06533_),
    .D(net843),
    .X(_06873_));
 mux2_1 _22763_ (.A0(net1375),
    .A1(\vmem[146] ),
    .S(_06873_),
    .X(_02005_));
 or4_1 _22764_ (.A(net747),
    .B(net629),
    .C(_06535_),
    .D(net845),
    .X(_06874_));
 mux2_1 _22765_ (.A0(net1379),
    .A1(\vmem[145] ),
    .S(_06874_),
    .X(_02006_));
 or4_1 _22766_ (.A(net727),
    .B(net612),
    .C(_06537_),
    .D(net827),
    .X(_06875_));
 mux2_1 _22767_ (.A0(net1341),
    .A1(\vmem[144] ),
    .S(_06875_),
    .X(_02007_));
 or4_1 _22768_ (.A(net736),
    .B(net618),
    .C(_06539_),
    .D(net836),
    .X(_06876_));
 mux2_1 _22769_ (.A0(net1358),
    .A1(\vmem[143] ),
    .S(_06876_),
    .X(_02008_));
 or4_1 _22770_ (.A(net741),
    .B(net622),
    .C(_06541_),
    .D(net839),
    .X(_06877_));
 mux2_1 _22771_ (.A0(net1368),
    .A1(\vmem[142] ),
    .S(_06877_),
    .X(_02009_));
 or4_1 _22772_ (.A(net739),
    .B(net621),
    .C(_06543_),
    .D(net840),
    .X(_06878_));
 mux2_1 _22773_ (.A0(net1365),
    .A1(\vmem[141] ),
    .S(_06878_),
    .X(_02010_));
 or4_1 _22774_ (.A(net753),
    .B(net634),
    .C(_06545_),
    .D(net850),
    .X(_06879_));
 mux2_1 _22775_ (.A0(net1386),
    .A1(\vmem[140] ),
    .S(_06879_),
    .X(_02011_));
 or4_1 _22776_ (.A(net738),
    .B(net618),
    .C(_06547_),
    .D(net837),
    .X(_06880_));
 mux2_1 _22777_ (.A0(net1358),
    .A1(\vmem[139] ),
    .S(_06880_),
    .X(_02012_));
 or4_1 _22778_ (.A(net730),
    .B(net614),
    .C(_06549_),
    .D(net830),
    .X(_06881_));
 mux2_1 _22779_ (.A0(net1345),
    .A1(\vmem[138] ),
    .S(_06881_),
    .X(_02013_));
 or4_1 _22780_ (.A(net728),
    .B(net612),
    .C(_06551_),
    .D(net828),
    .X(_06882_));
 mux2_1 _22781_ (.A0(net1342),
    .A1(\vmem[137] ),
    .S(_06882_),
    .X(_02014_));
 or4_1 _22782_ (.A(net724),
    .B(net609),
    .C(_06553_),
    .D(net824),
    .X(_06883_));
 mux2_1 _22783_ (.A0(net1335),
    .A1(\vmem[136] ),
    .S(_06883_),
    .X(_02015_));
 or4_1 _22784_ (.A(net733),
    .B(net617),
    .C(_06555_),
    .D(net833),
    .X(_06884_));
 mux2_1 _22785_ (.A0(net1351),
    .A1(\vmem[135] ),
    .S(_06884_),
    .X(_02016_));
 or4_1 _22786_ (.A(net754),
    .B(net637),
    .C(_06557_),
    .D(net849),
    .X(_06885_));
 mux2_1 _22787_ (.A0(net1386),
    .A1(\vmem[134] ),
    .S(_06885_),
    .X(_02017_));
 or4_1 _22788_ (.A(net726),
    .B(net605),
    .C(_06559_),
    .D(net825),
    .X(_06886_));
 mux2_1 _22789_ (.A0(net1336),
    .A1(\vmem[133] ),
    .S(_06886_),
    .X(_02018_));
 or4_1 _22790_ (.A(net750),
    .B(net632),
    .C(_06561_),
    .D(net847),
    .X(_06887_));
 mux2_1 _22791_ (.A0(net1383),
    .A1(\vmem[132] ),
    .S(_06887_),
    .X(_02019_));
 or4_1 _22792_ (.A(net720),
    .B(net608),
    .C(_06563_),
    .D(net821),
    .X(_06888_));
 mux2_1 _22793_ (.A0(net1328),
    .A1(\vmem[131] ),
    .S(_06888_),
    .X(_02020_));
 or4_1 _22794_ (.A(net744),
    .B(net626),
    .C(_06565_),
    .D(net843),
    .X(_06889_));
 mux2_1 _22795_ (.A0(net1354),
    .A1(\vmem[130] ),
    .S(_06889_),
    .X(_02021_));
 or4_1 _22796_ (.A(net746),
    .B(net627),
    .C(_06567_),
    .D(net845),
    .X(_06890_));
 mux2_1 _22797_ (.A0(net1377),
    .A1(\vmem[129] ),
    .S(_06890_),
    .X(_02022_));
 or4_1 _22798_ (.A(net723),
    .B(net607),
    .C(_06569_),
    .D(net823),
    .X(_06891_));
 mux2_1 _22799_ (.A0(net1341),
    .A1(\vmem[128] ),
    .S(_06891_),
    .X(_02023_));
 or4_1 _22800_ (.A(net772),
    .B(net650),
    .C(_06410_),
    .D(net832),
    .X(_06892_));
 mux2_1 _22801_ (.A0(net1347),
    .A1(\vmem[127] ),
    .S(_06892_),
    .X(_02024_));
 or4_1 _22802_ (.A(net782),
    .B(net659),
    .C(_06414_),
    .D(net839),
    .X(_06893_));
 mux2_1 _22803_ (.A0(net1367),
    .A1(\vmem[126] ),
    .S(_06893_),
    .X(_02025_));
 or4_1 _22804_ (.A(net781),
    .B(net661),
    .C(_06417_),
    .D(net838),
    .X(_06894_));
 mux2_1 _22805_ (.A0(net1352),
    .A1(\vmem[125] ),
    .S(_06894_),
    .X(_02026_));
 or4_1 _22806_ (.A(net790),
    .B(net666),
    .C(_06420_),
    .D(net844),
    .X(_06895_));
 mux2_1 _22807_ (.A0(net1378),
    .A1(\vmem[124] ),
    .S(_06895_),
    .X(_02027_));
 or4_1 _22808_ (.A(net779),
    .B(net657),
    .C(_06423_),
    .D(net835),
    .X(_06896_));
 mux2_1 _22809_ (.A0(net1360),
    .A1(\vmem[123] ),
    .S(_06896_),
    .X(_02028_));
 or4_1 _22810_ (.A(net770),
    .B(net649),
    .C(_06426_),
    .D(net830),
    .X(_06897_));
 mux2_1 _22811_ (.A0(net1346),
    .A1(\vmem[122] ),
    .S(_06897_),
    .X(_02029_));
 or4_1 _22812_ (.A(net786),
    .B(net664),
    .C(_06429_),
    .D(net842),
    .X(_06898_));
 mux2_1 _22813_ (.A0(net1371),
    .A1(\vmem[121] ),
    .S(_06898_),
    .X(_02030_));
 or4_1 _22814_ (.A(net763),
    .B(net644),
    .C(_06432_),
    .D(net825),
    .X(_06899_));
 mux2_1 _22815_ (.A0(net1337),
    .A1(\vmem[120] ),
    .S(_06899_),
    .X(_02031_));
 or4_1 _22816_ (.A(net775),
    .B(net652),
    .C(_06435_),
    .D(net833),
    .X(_06900_));
 mux2_1 _22817_ (.A0(net1351),
    .A1(\vmem[119] ),
    .S(_06900_),
    .X(_02032_));
 or4_1 _22818_ (.A(net798),
    .B(net673),
    .C(_06438_),
    .D(net849),
    .X(_06901_));
 mux2_1 _22819_ (.A0(net1392),
    .A1(\vmem[118] ),
    .S(_06901_),
    .X(_02033_));
 or4_1 _22820_ (.A(net759),
    .B(net640),
    .C(_06441_),
    .D(net821),
    .X(_06902_));
 mux2_1 _22821_ (.A0(net1329),
    .A1(\vmem[117] ),
    .S(_06902_),
    .X(_02034_));
 or4_1 _22822_ (.A(net794),
    .B(net668),
    .C(_06444_),
    .D(net848),
    .X(_06903_));
 mux2_1 _22823_ (.A0(net1384),
    .A1(\vmem[116] ),
    .S(_06903_),
    .X(_02035_));
 or4_1 _22824_ (.A(net759),
    .B(net640),
    .C(_06447_),
    .D(net821),
    .X(_06904_));
 mux2_1 _22825_ (.A0(net1329),
    .A1(\vmem[115] ),
    .S(_06904_),
    .X(_02036_));
 or4_1 _22826_ (.A(net792),
    .B(net670),
    .C(_06450_),
    .D(net846),
    .X(_06905_));
 mux2_1 _22827_ (.A0(net1380),
    .A1(\vmem[114] ),
    .S(_06905_),
    .X(_02037_));
 or4_1 _22828_ (.A(net786),
    .B(net664),
    .C(_06453_),
    .D(net842),
    .X(_06906_));
 mux2_1 _22829_ (.A0(net1372),
    .A1(\vmem[113] ),
    .S(_06906_),
    .X(_02038_));
 or4_1 _22830_ (.A(net766),
    .B(net646),
    .C(_06457_),
    .D(net827),
    .X(_06907_));
 mux2_1 _22831_ (.A0(net1341),
    .A1(\vmem[112] ),
    .S(_06907_),
    .X(_02039_));
 or4_1 _22832_ (.A(net772),
    .B(net650),
    .C(_06460_),
    .D(net832),
    .X(_06908_));
 mux2_1 _22833_ (.A0(net1347),
    .A1(\vmem[111] ),
    .S(_06908_),
    .X(_02040_));
 or4_1 _22834_ (.A(net782),
    .B(net659),
    .C(_06463_),
    .D(net839),
    .X(_06909_));
 mux2_1 _22835_ (.A0(net1367),
    .A1(\vmem[110] ),
    .S(_06909_),
    .X(_02041_));
 or4_1 _22836_ (.A(net781),
    .B(net661),
    .C(_06466_),
    .D(net838),
    .X(_06910_));
 mux2_1 _22837_ (.A0(net1364),
    .A1(\vmem[109] ),
    .S(_06910_),
    .X(_02042_));
 or4_1 _22838_ (.A(net790),
    .B(net667),
    .C(_06469_),
    .D(net845),
    .X(_06911_));
 mux2_1 _22839_ (.A0(net1377),
    .A1(\vmem[108] ),
    .S(_06911_),
    .X(_02043_));
 or4_1 _22840_ (.A(net779),
    .B(net657),
    .C(_06472_),
    .D(net835),
    .X(_06912_));
 mux2_1 _22841_ (.A0(net1360),
    .A1(\vmem[107] ),
    .S(_06912_),
    .X(_02044_));
 or4_1 _22842_ (.A(net770),
    .B(net649),
    .C(_06475_),
    .D(net830),
    .X(_06913_));
 mux2_1 _22843_ (.A0(net1345),
    .A1(\vmem[106] ),
    .S(_06913_),
    .X(_02045_));
 or4_1 _22844_ (.A(net786),
    .B(net664),
    .C(_06478_),
    .D(net842),
    .X(_06914_));
 mux2_1 _22845_ (.A0(net1371),
    .A1(\vmem[105] ),
    .S(_06914_),
    .X(_02046_));
 or4_1 _22846_ (.A(net765),
    .B(net643),
    .C(_06481_),
    .D(net826),
    .X(_06915_));
 mux2_1 _22847_ (.A0(net1338),
    .A1(\vmem[104] ),
    .S(_06915_),
    .X(_02047_));
 or4_1 _22848_ (.A(net775),
    .B(net652),
    .C(_06484_),
    .D(net833),
    .X(_06916_));
 mux2_1 _22849_ (.A0(net1351),
    .A1(\vmem[103] ),
    .S(_06916_),
    .X(_02048_));
 or4_1 _22850_ (.A(net798),
    .B(net673),
    .C(_06487_),
    .D(net849),
    .X(_06917_));
 mux2_1 _22851_ (.A0(net1392),
    .A1(\vmem[102] ),
    .S(_06917_),
    .X(_02049_));
 or4_1 _22852_ (.A(net759),
    .B(net640),
    .C(_06490_),
    .D(net821),
    .X(_06918_));
 mux2_1 _22853_ (.A0(net1329),
    .A1(\vmem[101] ),
    .S(_06918_),
    .X(_02050_));
 or4_1 _22854_ (.A(net794),
    .B(net668),
    .C(_06493_),
    .D(net848),
    .X(_06919_));
 mux2_1 _22855_ (.A0(net1384),
    .A1(\vmem[100] ),
    .S(_06919_),
    .X(_02051_));
 or4_1 _22856_ (.A(net758),
    .B(net640),
    .C(_06496_),
    .D(net820),
    .X(_06920_));
 mux2_1 _22857_ (.A0(net1327),
    .A1(\vmem[99] ),
    .S(_06920_),
    .X(_02052_));
 or4_1 _22858_ (.A(net792),
    .B(net670),
    .C(_06499_),
    .D(net846),
    .X(_06921_));
 mux2_1 _22859_ (.A0(net1380),
    .A1(\vmem[98] ),
    .S(_06921_),
    .X(_02053_));
 or4_1 _22860_ (.A(net791),
    .B(net667),
    .C(_06502_),
    .D(net845),
    .X(_06922_));
 mux2_1 _22861_ (.A0(net1379),
    .A1(\vmem[97] ),
    .S(_06922_),
    .X(_02054_));
 or4_1 _22862_ (.A(net766),
    .B(net645),
    .C(_06505_),
    .D(net827),
    .X(_06923_));
 mux2_1 _22863_ (.A0(net1341),
    .A1(\vmem[96] ),
    .S(_06923_),
    .X(_02055_));
 or4_1 _22864_ (.A(net772),
    .B(net651),
    .C(_06507_),
    .D(net832),
    .X(_06924_));
 mux2_1 _22865_ (.A0(net1348),
    .A1(\vmem[95] ),
    .S(_06924_),
    .X(_02056_));
 or4_1 _22866_ (.A(net782),
    .B(net659),
    .C(_06509_),
    .D(net839),
    .X(_06925_));
 mux2_1 _22867_ (.A0(net1367),
    .A1(\vmem[94] ),
    .S(_06925_),
    .X(_02057_));
 or4_1 _22868_ (.A(net774),
    .B(net653),
    .C(_06511_),
    .D(net834),
    .X(_06926_));
 mux2_1 _22869_ (.A0(net1354),
    .A1(\vmem[93] ),
    .S(_06926_),
    .X(_02058_));
 or4_1 _22870_ (.A(net799),
    .B(net671),
    .C(_06513_),
    .D(net850),
    .X(_06927_));
 mux2_1 _22871_ (.A0(net1387),
    .A1(\vmem[92] ),
    .S(_06927_),
    .X(_02059_));
 or4_1 _22872_ (.A(net777),
    .B(net655),
    .C(_06515_),
    .D(net835),
    .X(_06928_));
 mux2_1 _22873_ (.A0(net1357),
    .A1(\vmem[91] ),
    .S(_06928_),
    .X(_02060_));
 or4_1 _22874_ (.A(net770),
    .B(net649),
    .C(_06517_),
    .D(net831),
    .X(_06929_));
 mux2_1 _22875_ (.A0(net1346),
    .A1(\vmem[90] ),
    .S(_06929_),
    .X(_02061_));
 or4_1 _22876_ (.A(net769),
    .B(net648),
    .C(_06519_),
    .D(net829),
    .X(_06930_));
 mux2_1 _22877_ (.A0(net1344),
    .A1(\vmem[89] ),
    .S(_06930_),
    .X(_02062_));
 or4_1 _22878_ (.A(net765),
    .B(net643),
    .C(_06521_),
    .D(net826),
    .X(_06931_));
 mux2_1 _22879_ (.A0(net1338),
    .A1(\vmem[88] ),
    .S(_06931_),
    .X(_02063_));
 or4_1 _22880_ (.A(net771),
    .B(net649),
    .C(_06523_),
    .D(net831),
    .X(_06932_));
 mux2_1 _22881_ (.A0(net1346),
    .A1(\vmem[87] ),
    .S(_06932_),
    .X(_02064_));
 or4_1 _22882_ (.A(net798),
    .B(net672),
    .C(_06525_),
    .D(net849),
    .X(_06933_));
 mux2_1 _22883_ (.A0(net1391),
    .A1(\vmem[86] ),
    .S(_06933_),
    .X(_02065_));
 or4_1 _22884_ (.A(net760),
    .B(net642),
    .C(_06527_),
    .D(net822),
    .X(_06934_));
 mux2_1 _22885_ (.A0(net1331),
    .A1(\vmem[85] ),
    .S(_06934_),
    .X(_02066_));
 or4_1 _22886_ (.A(net793),
    .B(net669),
    .C(_06529_),
    .D(net847),
    .X(_06935_));
 mux2_1 _22887_ (.A0(net1383),
    .A1(\vmem[84] ),
    .S(_06935_),
    .X(_02067_));
 or4_1 _22888_ (.A(net758),
    .B(net640),
    .C(_06531_),
    .D(net820),
    .X(_06936_));
 mux2_1 _22889_ (.A0(net1327),
    .A1(\vmem[83] ),
    .S(_06936_),
    .X(_02068_));
 or4_1 _22890_ (.A(net792),
    .B(net670),
    .C(_06533_),
    .D(net846),
    .X(_06937_));
 mux2_1 _22891_ (.A0(net1382),
    .A1(\vmem[82] ),
    .S(_06937_),
    .X(_02069_));
 or4_1 _22892_ (.A(net786),
    .B(net664),
    .C(_06535_),
    .D(net842),
    .X(_06938_));
 mux2_1 _22893_ (.A0(net1372),
    .A1(\vmem[81] ),
    .S(_06938_),
    .X(_02070_));
 or4_1 _22894_ (.A(net766),
    .B(net645),
    .C(_06537_),
    .D(net827),
    .X(_06939_));
 mux2_1 _22895_ (.A0(net1340),
    .A1(\vmem[80] ),
    .S(_06939_),
    .X(_02071_));
 or4_1 _22896_ (.A(net777),
    .B(net655),
    .C(_06539_),
    .D(net836),
    .X(_06940_));
 mux2_1 _22897_ (.A0(net1348),
    .A1(\vmem[79] ),
    .S(_06940_),
    .X(_02072_));
 or4_1 _22898_ (.A(net782),
    .B(net659),
    .C(_06541_),
    .D(net839),
    .X(_06941_));
 mux2_1 _22899_ (.A0(net1364),
    .A1(\vmem[78] ),
    .S(_06941_),
    .X(_02073_));
 or4_1 _22900_ (.A(net778),
    .B(net656),
    .C(_06543_),
    .D(net836),
    .X(_06942_));
 mux2_1 _22901_ (.A0(net1358),
    .A1(\vmem[77] ),
    .S(_06942_),
    .X(_02074_));
 or4_1 _22902_ (.A(net796),
    .B(net671),
    .C(_06545_),
    .D(net850),
    .X(_06943_));
 mux2_1 _22903_ (.A0(net1387),
    .A1(\vmem[76] ),
    .S(_06943_),
    .X(_02075_));
 or4_1 _22904_ (.A(net779),
    .B(net657),
    .C(_06547_),
    .D(net835),
    .X(_06944_));
 mux2_1 _22905_ (.A0(net1357),
    .A1(\vmem[75] ),
    .S(_06944_),
    .X(_02076_));
 or4_1 _22906_ (.A(net770),
    .B(net649),
    .C(_06549_),
    .D(net830),
    .X(_06945_));
 mux2_1 _22907_ (.A0(net1345),
    .A1(\vmem[74] ),
    .S(_06945_),
    .X(_02077_));
 or4_1 _22908_ (.A(net769),
    .B(net648),
    .C(_06551_),
    .D(net829),
    .X(_06946_));
 mux2_1 _22909_ (.A0(net1344),
    .A1(\vmem[73] ),
    .S(_06946_),
    .X(_02078_));
 or4_1 _22910_ (.A(net763),
    .B(net644),
    .C(_06553_),
    .D(net824),
    .X(_06947_));
 mux2_1 _22911_ (.A0(net1335),
    .A1(\vmem[72] ),
    .S(_06947_),
    .X(_02079_));
 or4_1 _22912_ (.A(net771),
    .B(net649),
    .C(_06555_),
    .D(net831),
    .X(_06948_));
 mux2_1 _22913_ (.A0(net1346),
    .A1(\vmem[71] ),
    .S(_06948_),
    .X(_02080_));
 or4_1 _22914_ (.A(net798),
    .B(net672),
    .C(_06557_),
    .D(net849),
    .X(_06949_));
 mux2_1 _22915_ (.A0(net1392),
    .A1(\vmem[70] ),
    .S(_06949_),
    .X(_02081_));
 or4_1 _22916_ (.A(net761),
    .B(net641),
    .C(_06559_),
    .D(net822),
    .X(_06950_));
 mux2_1 _22917_ (.A0(net1331),
    .A1(\vmem[69] ),
    .S(_06950_),
    .X(_02082_));
 or4_1 _22918_ (.A(net794),
    .B(net668),
    .C(_06561_),
    .D(net848),
    .X(_06951_));
 mux2_1 _22919_ (.A0(net1384),
    .A1(\vmem[68] ),
    .S(_06951_),
    .X(_02083_));
 or4_1 _22920_ (.A(net759),
    .B(net642),
    .C(_06563_),
    .D(net822),
    .X(_06952_));
 mux2_1 _22921_ (.A0(net1329),
    .A1(\vmem[67] ),
    .S(_06952_),
    .X(_02084_));
 or4_1 _22922_ (.A(net792),
    .B(net670),
    .C(_06565_),
    .D(net846),
    .X(_06953_));
 mux2_1 _22923_ (.A0(net1380),
    .A1(\vmem[66] ),
    .S(_06953_),
    .X(_02085_));
 or4_1 _22924_ (.A(net789),
    .B(net666),
    .C(_06567_),
    .D(net844),
    .X(_06954_));
 mux2_1 _22925_ (.A0(net1379),
    .A1(\vmem[65] ),
    .S(_06954_),
    .X(_02086_));
 or4_1 _22926_ (.A(net766),
    .B(net645),
    .C(_06569_),
    .D(net827),
    .X(_06955_));
 mux2_1 _22927_ (.A0(net1340),
    .A1(\vmem[64] ),
    .S(_06955_),
    .X(_02087_));
 or4_1 _22928_ (.A(net735),
    .B(net655),
    .C(_06410_),
    .D(net836),
    .X(_06956_));
 mux2_1 _22929_ (.A0(net1356),
    .A1(\vmem[63] ),
    .S(_06956_),
    .X(_02088_));
 or4_1 _22930_ (.A(net741),
    .B(net660),
    .C(_06414_),
    .D(net840),
    .X(_06957_));
 mux2_1 _22931_ (.A0(net1368),
    .A1(\vmem[62] ),
    .S(_06957_),
    .X(_02089_));
 or4_1 _22932_ (.A(net739),
    .B(net661),
    .C(_06417_),
    .D(net838),
    .X(_06958_));
 mux2_1 _22933_ (.A0(net1364),
    .A1(\vmem[61] ),
    .S(_06958_),
    .X(_02090_));
 or4_1 _22934_ (.A(net747),
    .B(net666),
    .C(_06420_),
    .D(net845),
    .X(_06959_));
 mux2_1 _22935_ (.A0(net1377),
    .A1(\vmem[60] ),
    .S(_06959_),
    .X(_02091_));
 or4_1 _22936_ (.A(net737),
    .B(net657),
    .C(_06423_),
    .D(net835),
    .X(_06960_));
 mux2_1 _22937_ (.A0(net1360),
    .A1(\vmem[59] ),
    .S(_06960_),
    .X(_02092_));
 or4_1 _22938_ (.A(net730),
    .B(net654),
    .C(_06426_),
    .D(net831),
    .X(_06961_));
 mux2_1 _22939_ (.A0(net1350),
    .A1(\vmem[58] ),
    .S(_06961_),
    .X(_02093_));
 or4_1 _22940_ (.A(net743),
    .B(net664),
    .C(_06429_),
    .D(net842),
    .X(_06962_));
 mux2_1 _22941_ (.A0(net1371),
    .A1(\vmem[57] ),
    .S(_06962_),
    .X(_02094_));
 or4_1 _22942_ (.A(net725),
    .B(net643),
    .C(_06432_),
    .D(net826),
    .X(_06963_));
 mux2_1 _22943_ (.A0(net1338),
    .A1(\vmem[56] ),
    .S(_06963_),
    .X(_02095_));
 or4_1 _22944_ (.A(net733),
    .B(net652),
    .C(_06435_),
    .D(net833),
    .X(_06964_));
 mux2_1 _22945_ (.A0(net1351),
    .A1(\vmem[55] ),
    .S(_06964_),
    .X(_02096_));
 or4_1 _22946_ (.A(net754),
    .B(net672),
    .C(_06438_),
    .D(net851),
    .X(_06965_));
 mux2_1 _22947_ (.A0(net1391),
    .A1(\vmem[54] ),
    .S(_06965_),
    .X(_02097_));
 or4_1 _22948_ (.A(net720),
    .B(net640),
    .C(_06441_),
    .D(net821),
    .X(_06966_));
 mux2_1 _22949_ (.A0(net1329),
    .A1(\vmem[53] ),
    .S(_06966_),
    .X(_02098_));
 or4_1 _22950_ (.A(net749),
    .B(net670),
    .C(_06444_),
    .D(net851),
    .X(_06967_));
 mux2_1 _22951_ (.A0(net1382),
    .A1(\vmem[52] ),
    .S(_06967_),
    .X(_02099_));
 or4_1 _22952_ (.A(net720),
    .B(net640),
    .C(_06447_),
    .D(net821),
    .X(_06968_));
 mux2_1 _22953_ (.A0(net1329),
    .A1(\vmem[51] ),
    .S(_06968_),
    .X(_02100_));
 or4_1 _22954_ (.A(net749),
    .B(net670),
    .C(_06450_),
    .D(net846),
    .X(_06969_));
 mux2_1 _22955_ (.A0(net1380),
    .A1(\vmem[50] ),
    .S(_06969_),
    .X(_02101_));
 or4_1 _22956_ (.A(net743),
    .B(net664),
    .C(_06453_),
    .D(net843),
    .X(_06970_));
 mux2_1 _22957_ (.A0(net1372),
    .A1(\vmem[49] ),
    .S(_06970_),
    .X(_02102_));
 or4_1 _22958_ (.A(net727),
    .B(net645),
    .C(_06457_),
    .D(net827),
    .X(_06971_));
 mux2_1 _22959_ (.A0(net1340),
    .A1(\vmem[48] ),
    .S(_06971_),
    .X(_02103_));
 or4_1 _22960_ (.A(net731),
    .B(net650),
    .C(_06460_),
    .D(net832),
    .X(_06972_));
 mux2_1 _22961_ (.A0(net1348),
    .A1(\vmem[47] ),
    .S(_06972_),
    .X(_02104_));
 or4_1 _22962_ (.A(net750),
    .B(net669),
    .C(_06463_),
    .D(net847),
    .X(_06973_));
 mux2_1 _22963_ (.A0(net1383),
    .A1(\vmem[46] ),
    .S(_06973_),
    .X(_02105_));
 or4_1 _22964_ (.A(net739),
    .B(net661),
    .C(_06466_),
    .D(net838),
    .X(_06974_));
 mux2_1 _22965_ (.A0(net1365),
    .A1(\vmem[45] ),
    .S(_06974_),
    .X(_02106_));
 or4_1 _22966_ (.A(net747),
    .B(net666),
    .C(_06469_),
    .D(net844),
    .X(_06975_));
 mux2_1 _22967_ (.A0(net1378),
    .A1(\vmem[44] ),
    .S(_06975_),
    .X(_02107_));
 or4_1 _22968_ (.A(net737),
    .B(net658),
    .C(_06472_),
    .D(net835),
    .X(_06976_));
 mux2_1 _22969_ (.A0(net1360),
    .A1(\vmem[43] ),
    .S(_06976_),
    .X(_02108_));
 or4_1 _22970_ (.A(net730),
    .B(net649),
    .C(_06475_),
    .D(net830),
    .X(_06977_));
 mux2_1 _22971_ (.A0(net1346),
    .A1(\vmem[42] ),
    .S(_06977_),
    .X(_02109_));
 or4_1 _22972_ (.A(net743),
    .B(net664),
    .C(_06478_),
    .D(net842),
    .X(_06978_));
 mux2_1 _22973_ (.A0(net1371),
    .A1(\vmem[41] ),
    .S(_06978_),
    .X(_02110_));
 or4_1 _22974_ (.A(net725),
    .B(net643),
    .C(_06481_),
    .D(net826),
    .X(_06979_));
 mux2_1 _22975_ (.A0(net1338),
    .A1(\vmem[40] ),
    .S(_06979_),
    .X(_02111_));
 or4_1 _22976_ (.A(net733),
    .B(net652),
    .C(_06484_),
    .D(net833),
    .X(_06980_));
 mux2_1 _22977_ (.A0(net1351),
    .A1(\vmem[39] ),
    .S(_06980_),
    .X(_02112_));
 or4_1 _22978_ (.A(net754),
    .B(net673),
    .C(_06487_),
    .D(net851),
    .X(_06981_));
 mux2_1 _22979_ (.A0(net1391),
    .A1(\vmem[38] ),
    .S(_06981_),
    .X(_02113_));
 or4_1 _22980_ (.A(net720),
    .B(net642),
    .C(_06490_),
    .D(net821),
    .X(_06982_));
 mux2_1 _22981_ (.A0(net1329),
    .A1(\vmem[37] ),
    .S(_06982_),
    .X(_02114_));
 or4_1 _22982_ (.A(net749),
    .B(net670),
    .C(_06493_),
    .D(net851),
    .X(_06983_));
 mux2_1 _22983_ (.A0(net1382),
    .A1(\vmem[36] ),
    .S(_06983_),
    .X(_02115_));
 or4_1 _22984_ (.A(net720),
    .B(net640),
    .C(_06496_),
    .D(net821),
    .X(_06984_));
 mux2_1 _22985_ (.A0(net1328),
    .A1(\vmem[35] ),
    .S(_06984_),
    .X(_02116_));
 or4_1 _22986_ (.A(net749),
    .B(net670),
    .C(_06499_),
    .D(net846),
    .X(_06985_));
 mux2_1 _22987_ (.A0(net1380),
    .A1(\vmem[34] ),
    .S(_06985_),
    .X(_02117_));
 or4_1 _22988_ (.A(net748),
    .B(net667),
    .C(_06502_),
    .D(net845),
    .X(_06986_));
 mux2_1 _22989_ (.A0(net1372),
    .A1(\vmem[33] ),
    .S(_06986_),
    .X(_02118_));
 or4_1 _22990_ (.A(net727),
    .B(net645),
    .C(_06505_),
    .D(net827),
    .X(_06987_));
 mux2_1 _22991_ (.A0(net1340),
    .A1(\vmem[32] ),
    .S(_06987_),
    .X(_02119_));
 or4_1 _22992_ (.A(net731),
    .B(net655),
    .C(_06507_),
    .D(net836),
    .X(_06988_));
 mux2_1 _22993_ (.A0(net1347),
    .A1(\vmem[31] ),
    .S(_06988_),
    .X(_02120_));
 or4_1 _22994_ (.A(net740),
    .B(net659),
    .C(_06509_),
    .D(net839),
    .X(_06989_));
 mux2_1 _22995_ (.A0(net1367),
    .A1(\vmem[30] ),
    .S(_06989_),
    .X(_02121_));
 or4_1 _22996_ (.A(net734),
    .B(net653),
    .C(_06511_),
    .D(net834),
    .X(_06990_));
 mux2_1 _22997_ (.A0(net1352),
    .A1(\vmem[29] ),
    .S(_06990_),
    .X(_02122_));
 or4_1 _22998_ (.A(net756),
    .B(net671),
    .C(_06513_),
    .D(net850),
    .X(_06991_));
 mux2_1 _22999_ (.A0(net1387),
    .A1(\vmem[28] ),
    .S(_06991_),
    .X(_02123_));
 or4_1 _23000_ (.A(net737),
    .B(net657),
    .C(_06515_),
    .D(net835),
    .X(_06992_));
 mux2_1 _23001_ (.A0(net1360),
    .A1(\vmem[27] ),
    .S(_06992_),
    .X(_02124_));
 or4_1 _23002_ (.A(net730),
    .B(net649),
    .C(_06517_),
    .D(net830),
    .X(_06993_));
 mux2_1 _23003_ (.A0(net1346),
    .A1(\vmem[26] ),
    .S(_06993_),
    .X(_02125_));
 or4_1 _23004_ (.A(_03766_),
    .B(net648),
    .C(_06519_),
    .D(net829),
    .X(_06994_));
 mux2_1 _23005_ (.A0(net1344),
    .A1(\vmem[25] ),
    .S(_06994_),
    .X(_02126_));
 or4_1 _23006_ (.A(net725),
    .B(net643),
    .C(_06521_),
    .D(net826),
    .X(_06995_));
 mux2_1 _23007_ (.A0(net1338),
    .A1(\vmem[24] ),
    .S(_06995_),
    .X(_02127_));
 or4_1 _23008_ (.A(net730),
    .B(net654),
    .C(_06523_),
    .D(net831),
    .X(_06996_));
 mux2_1 _23009_ (.A0(net1350),
    .A1(\vmem[23] ),
    .S(_06996_),
    .X(_02128_));
 or4_1 _23010_ (.A(net755),
    .B(net673),
    .C(_06525_),
    .D(net850),
    .X(_06997_));
 mux2_1 _23011_ (.A0(net1391),
    .A1(\vmem[22] ),
    .S(_06997_),
    .X(_02129_));
 or4_1 _23012_ (.A(net722),
    .B(net641),
    .C(_06527_),
    .D(net822),
    .X(_06998_));
 mux2_1 _23013_ (.A0(net1331),
    .A1(\vmem[21] ),
    .S(_06998_),
    .X(_02130_));
 or4_1 _23014_ (.A(net750),
    .B(net668),
    .C(_06529_),
    .D(net848),
    .X(_06999_));
 mux2_1 _23015_ (.A0(net1384),
    .A1(\vmem[20] ),
    .S(_06999_),
    .X(_02131_));
 or4_1 _23016_ (.A(net720),
    .B(net640),
    .C(_06531_),
    .D(net820),
    .X(_07000_));
 mux2_1 _23017_ (.A0(net1327),
    .A1(\vmem[19] ),
    .S(_07000_),
    .X(_02132_));
 or4_1 _23018_ (.A(net749),
    .B(net670),
    .C(_06533_),
    .D(net846),
    .X(_07001_));
 mux2_1 _23019_ (.A0(net1380),
    .A1(\vmem[18] ),
    .S(_07001_),
    .X(_02133_));
 or4_1 _23020_ (.A(net745),
    .B(net665),
    .C(_06535_),
    .D(net852),
    .X(_07002_));
 mux2_1 _23021_ (.A0(net1374),
    .A1(\vmem[17] ),
    .S(_07002_),
    .X(_02134_));
 or4_1 _23022_ (.A(net724),
    .B(net644),
    .C(_06537_),
    .D(net825),
    .X(_07003_));
 mux2_1 _23023_ (.A0(net1336),
    .A1(\vmem[16] ),
    .S(_07003_),
    .X(_02135_));
 or4_1 _23024_ (.A(net735),
    .B(net655),
    .C(_06539_),
    .D(net836),
    .X(_07004_));
 mux2_1 _23025_ (.A0(net1356),
    .A1(\vmem[15] ),
    .S(_07004_),
    .X(_02136_));
 or4_1 _23026_ (.A(net740),
    .B(net659),
    .C(_06541_),
    .D(net839),
    .X(_07005_));
 mux2_1 _23027_ (.A0(net1367),
    .A1(\vmem[14] ),
    .S(_07005_),
    .X(_02137_));
 or4_1 _23028_ (.A(net734),
    .B(net653),
    .C(_06543_),
    .D(net834),
    .X(_07006_));
 mux2_1 _23029_ (.A0(net1352),
    .A1(\vmem[13] ),
    .S(_07006_),
    .X(_02138_));
 or4_1 _23030_ (.A(net756),
    .B(net671),
    .C(_06545_),
    .D(net850),
    .X(_07007_));
 mux2_1 _23031_ (.A0(net1387),
    .A1(\vmem[12] ),
    .S(_07007_),
    .X(_02139_));
 or4_1 _23032_ (.A(net737),
    .B(net657),
    .C(_06547_),
    .D(net835),
    .X(_07008_));
 mux2_1 _23033_ (.A0(net1360),
    .A1(\vmem[11] ),
    .S(_07008_),
    .X(_02140_));
 or4_1 _23034_ (.A(net730),
    .B(net649),
    .C(_06549_),
    .D(net830),
    .X(_07009_));
 mux2_1 _23035_ (.A0(net1345),
    .A1(\vmem[10] ),
    .S(_07009_),
    .X(_02141_));
 or4_1 _23036_ (.A(_03766_),
    .B(net648),
    .C(_06551_),
    .D(net829),
    .X(_07010_));
 mux2_1 _23037_ (.A0(net1344),
    .A1(\vmem[9] ),
    .S(_07010_),
    .X(_02142_));
 or4_1 _23038_ (.A(net725),
    .B(net643),
    .C(_06553_),
    .D(net826),
    .X(_07011_));
 mux2_1 _23039_ (.A0(net1338),
    .A1(\vmem[8] ),
    .S(_07011_),
    .X(_02143_));
 or4_1 _23040_ (.A(net732),
    .B(net649),
    .C(_06555_),
    .D(net831),
    .X(_07012_));
 mux2_1 _23041_ (.A0(net1350),
    .A1(\vmem[7] ),
    .S(_07012_),
    .X(_02144_));
 or4_1 _23042_ (.A(net755),
    .B(net673),
    .C(_06557_),
    .D(net850),
    .X(_07013_));
 mux2_1 _23043_ (.A0(net1391),
    .A1(\vmem[6] ),
    .S(_07013_),
    .X(_02145_));
 or4_1 _23044_ (.A(net721),
    .B(net641),
    .C(_06559_),
    .D(net822),
    .X(_07014_));
 mux2_1 _23045_ (.A0(net1331),
    .A1(\vmem[5] ),
    .S(_07014_),
    .X(_02146_));
 or4_1 _23046_ (.A(net751),
    .B(net668),
    .C(_06561_),
    .D(net848),
    .X(_07015_));
 mux2_1 _23047_ (.A0(net1384),
    .A1(\vmem[4] ),
    .S(_07015_),
    .X(_02147_));
 or4_1 _23048_ (.A(net720),
    .B(net642),
    .C(_06563_),
    .D(net820),
    .X(_07016_));
 mux2_1 _23049_ (.A0(net1329),
    .A1(\vmem[3] ),
    .S(_07016_),
    .X(_02148_));
 or4_1 _23050_ (.A(net749),
    .B(net670),
    .C(_06565_),
    .D(net846),
    .X(_07017_));
 mux2_1 _23051_ (.A0(net1382),
    .A1(\vmem[2] ),
    .S(_07017_),
    .X(_02149_));
 or4_1 _23052_ (.A(net745),
    .B(net665),
    .C(_06567_),
    .D(net852),
    .X(_07018_));
 mux2_1 _23053_ (.A0(net1374),
    .A1(\vmem[1] ),
    .S(_07018_),
    .X(_02150_));
 or4_1 _23054_ (.A(net727),
    .B(net645),
    .C(_06569_),
    .D(net827),
    .X(_07019_));
 mux2_1 _23055_ (.A0(net1340),
    .A1(\vmem[0] ),
    .S(_07019_),
    .X(_02151_));
 nand2_1 _23056_ (.A(net1398),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_i ),
    .Y(_00259_));
 or2_1 _23057_ (.A(net1446),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_i ),
    .X(_00258_));
 nand2_1 _23058_ (.A(net1398),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.sl_i ),
    .Y(_00253_));
 or2_1 _23059_ (.A(net1452),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.sl_i ),
    .X(_00252_));
 or2_1 _23060_ (.A(net1452),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ),
    .X(_00250_));
 nand2_1 _23061_ (.A(net1398),
    .B(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ),
    .Y(_00249_));
 inv_2 _23062_ (.A(_00206_),
    .Y(\digitop_pav2.sync_inst.inst_clkx.en_blf_fc_b ));
 or2_1 _23063_ (.A(net1273),
    .B(_00267_),
    .X(\digitop_pav2.sync_inst.inst_clkx.g_invent ));
 inv_2 _23064_ (.A(net1697),
    .Y(_00171_));
 inv_2 _23065_ (.A(net1213),
    .Y(_00172_));
 inv_2 _23066_ (.A(net1213),
    .Y(_00173_));
 inv_2 _23067_ (.A(net1204),
    .Y(_00174_));
 inv_2 _23068_ (.A(net1201),
    .Y(_00175_));
 inv_2 _23069_ (.A(net1201),
    .Y(_00176_));
 inv_2 _23070_ (.A(net1207),
    .Y(_00177_));
 inv_2 _23071_ (.A(net1205),
    .Y(_00178_));
 inv_2 _23072_ (.A(net1206),
    .Y(_00179_));
 inv_2 _23073_ (.A(net1206),
    .Y(_00180_));
 inv_2 _23074_ (.A(net1204),
    .Y(_00181_));
 inv_2 _23075_ (.A(net1203),
    .Y(_00182_));
 inv_2 _23076_ (.A(net1206),
    .Y(_00183_));
 inv_2 _23077_ (.A(net1201),
    .Y(_00184_));
 inv_2 _23078_ (.A(net1207),
    .Y(_00185_));
 inv_2 _23079_ (.A(net1206),
    .Y(_00186_));
 inv_2 _23080_ (.A(net1204),
    .Y(_00187_));
 inv_2 _23081_ (.A(net1202),
    .Y(_00188_));
 inv_2 _23082_ (.A(net1210),
    .Y(_00189_));
 inv_2 _23083_ (.A(net1211),
    .Y(_00190_));
 inv_2 _23084_ (.A(net1205),
    .Y(_00191_));
 inv_2 _23085_ (.A(net1208),
    .Y(_00192_));
 inv_2 _23086_ (.A(net1202),
    .Y(_00193_));
 inv_2 _23087_ (.A(net1209),
    .Y(_00194_));
 inv_2 _23088_ (.A(net1204),
    .Y(_00195_));
 inv_2 _23089_ (.A(net1204),
    .Y(_00196_));
 inv_2 _23090_ (.A(net1211),
    .Y(_00197_));
 inv_2 _23091_ (.A(net1205),
    .Y(_00198_));
 inv_2 _23092_ (.A(net1205),
    .Y(_00199_));
 inv_2 _23093_ (.A(net1207),
    .Y(_00200_));
 inv_2 _23094_ (.A(net1204),
    .Y(_00201_));
 inv_2 _23095_ (.A(net1205),
    .Y(_00202_));
 nand2_1 _23096_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.dis_blf_fc_b ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.en_blf_fc_b ),
    .Y(_00209_));
 nand2_2 _23097_ (.A(net1725),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.en_blf_fc_b ),
    .Y(_00210_));
 nand2_1 _23098_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.dis_blf_fc_b ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.en_blf_fc_b ),
    .Y(_00211_));
 clkbuf_1 _23099_ (.A(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_en.slow_clk_en_b_ff2_i ),
    .X(_00580_));
 nor2_1 _23100_ (.A(net1397),
    .B(net156),
    .Y(_00217_));
 nor2_1 _23101_ (.A(net1397),
    .B(net156),
    .Y(_00218_));
 nor2_1 _23102_ (.A(net1397),
    .B(net156),
    .Y(_00219_));
 nor2_1 _23103_ (.A(net1396),
    .B(net156),
    .Y(_00220_));
 nor2_1 _23104_ (.A(net1396),
    .B(net156),
    .Y(_00221_));
 nor2_1 _23105_ (.A(net1399),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.fm0x_mod_en_i ),
    .Y(_00222_));
 nor2_1 _23106_ (.A(net1399),
    .B(\digitop_pav2.proc_ctrl_inst.cmdfsm.fm0x_mod_en_i ),
    .Y(_00223_));
 nor2_1 _23107_ (.A(net1396),
    .B(net967),
    .Y(_00225_));
 nor2_1 _23108_ (.A(net1396),
    .B(net968),
    .Y(_00226_));
 nor2_1 _23109_ (.A(net1397),
    .B(net967),
    .Y(_00227_));
 nor2_1 _23110_ (.A(net1397),
    .B(net967),
    .Y(_00228_));
 nor2_1 _23111_ (.A(net1397),
    .B(net967),
    .Y(_00229_));
 nor2_1 _23112_ (.A(net1397),
    .B(net967),
    .Y(_00230_));
 nor2_1 _23113_ (.A(net1397),
    .B(net967),
    .Y(_00231_));
 nor2_1 _23114_ (.A(net1396),
    .B(net967),
    .Y(_00232_));
 nor2_1 _23115_ (.A(net1396),
    .B(net967),
    .Y(_00233_));
 nor2_1 _23116_ (.A(net1396),
    .B(net967),
    .Y(_00234_));
 nor2_1 _23117_ (.A(net1396),
    .B(net967),
    .Y(_00235_));
 nor2_1 _23118_ (.A(net1396),
    .B(net968),
    .Y(_00236_));
 inv_2 _23119_ (.A(\digitop_pav2.pie_inst.fsm.clk_i ),
    .Y(_00238_));
 inv_2 _23120_ (.A(\digitop_pav2.pie_inst.fsm.clk_i ),
    .Y(_00239_));
 inv_2 _23121_ (.A(\digitop_pav2.pie_inst.fsm.clk_i ),
    .Y(_00240_));
 inv_2 _23122_ (.A(\digitop_pav2.pie_inst.fsm.clk_i ),
    .Y(_00241_));
 inv_2 _23123_ (.A(\digitop_pav2.pie_inst.fsm.clk_i ),
    .Y(_00242_));
 inv_2 _23124_ (.A(\digitop_pav2.pie_inst.fsm.clk_i ),
    .Y(_00243_));
 inv_2 _23125_ (.A(\digitop_pav2.pie_inst.fsm.clk_i ),
    .Y(_00244_));
 inv_2 _23126_ (.A(\digitop_pav2.pie_inst.fsm.clk_i ),
    .Y(_00245_));
 clkbuf_1 _23127_ (.A(\digitop_pav2.pie_inst.fsm.comp_delimiter_ff ),
    .X(_01046_));
 inv_2 _23128_ (.A(\digitop_pav2.clkx_invent_clk ),
    .Y(_00251_));
 inv_2 _23129_ (.A(\digitop_pav2.clkx_invent_clk ),
    .Y(_00254_));
 inv_2 _23130_ (.A(\digitop_pav2.clkx_invent_clk ),
    .Y(_00257_));
 inv_2 _23131_ (.A(\digitop_pav2.clkx_invent_clk ),
    .Y(_00260_));
 inv_2 _23132_ (.A(\digitop_pav2.clkx_invent_clk ),
    .Y(_00263_));
 inv_2 _23133_ (.A(\digitop_pav2.clkx_invent_clk ),
    .Y(_00266_));
 or4_1 _23134_ (.A(net1678),
    .B(net1277),
    .C(net1669),
    .D(net1675),
    .X(_00268_));
 or4_1 _23135_ (.A(net1274),
    .B(net1672),
    .C(net1279),
    .D(net1282),
    .X(_00269_));
 or4_1 _23136_ (.A(net1274),
    .B(net1672),
    .C(net1669),
    .D(net1282),
    .X(_00270_));
 or4_1 _23137_ (.A(net1678),
    .B(net1277),
    .C(net1669),
    .D(net1675),
    .X(_00271_));
 or4_1 _23138_ (.A(net1274),
    .B(net1672),
    .C(net1279),
    .D(net1282),
    .X(_00272_));
 or4_1 _23139_ (.A(net1274),
    .B(net1672),
    .C(net1279),
    .D(net1282),
    .X(_00273_));
 or4_1 _23140_ (.A(net1678),
    .B(net1672),
    .C(net1279),
    .D(net1282),
    .X(_00274_));
 or4_1 _23141_ (.A(net1274),
    .B(net1277),
    .C(net1669),
    .D(net1282),
    .X(_00275_));
 or4_1 _23142_ (.A(net1678),
    .B(net1672),
    .C(net1279),
    .D(net1282),
    .X(_00276_));
 and2_1 _23143_ (.A(net1438),
    .B(net1220),
    .X(_00278_));
 and2_1 _23144_ (.A(net1438),
    .B(net1221),
    .X(_00279_));
 and2_1 _23145_ (.A(net1438),
    .B(net1222),
    .X(_00280_));
 and2_1 _23146_ (.A(net1438),
    .B(net1222),
    .X(_00281_));
 and2_1 _23147_ (.A(net1443),
    .B(net1221),
    .X(_00282_));
 and2_1 _23148_ (.A(net1438),
    .B(net1222),
    .X(_00283_));
 and2_1 _23149_ (.A(net1438),
    .B(net1220),
    .X(_00284_));
 and2_1 _23150_ (.A(net1440),
    .B(net1220),
    .X(_00285_));
 and2_1 _23151_ (.A(net1440),
    .B(net1220),
    .X(_00286_));
 and2_1 _23152_ (.A(net1440),
    .B(net1222),
    .X(_00287_));
 and2_1 _23153_ (.A(net1440),
    .B(net1222),
    .X(_00288_));
 and2_1 _23154_ (.A(net1440),
    .B(net1222),
    .X(_00289_));
 and2_1 _23155_ (.A(net1443),
    .B(net1220),
    .X(_00290_));
 and2_1 _23156_ (.A(net1440),
    .B(net1220),
    .X(_00291_));
 and2_1 _23157_ (.A(net1440),
    .B(net1220),
    .X(_00292_));
 inv_2 _23158_ (.A(\digitop_pav2.clkx_fm0x_clk ),
    .Y(_00294_));
 and2_1 _23159_ (.A(net1440),
    .B(net1220),
    .X(_00295_));
 and2_1 _23160_ (.A(net1440),
    .B(net1220),
    .X(_00296_));
 and2_1 _23161_ (.A(net1438),
    .B(net1221),
    .X(_00297_));
 and2_1 _23162_ (.A(net1438),
    .B(net1220),
    .X(_00298_));
 and2_1 _23163_ (.A(net1439),
    .B(net1221),
    .X(_00299_));
 and2_1 _23164_ (.A(net1439),
    .B(net1221),
    .X(_00300_));
 and2_1 _23165_ (.A(net1439),
    .B(net1221),
    .X(_00301_));
 and2_1 _23166_ (.A(net1438),
    .B(net1221),
    .X(_00302_));
 and2_1 _23167_ (.A(net1439),
    .B(net1221),
    .X(_00303_));
 clkbuf_1 _23168_ (.A(net1302),
    .X(_01194_));
 inv_2 _23169_ (.A(net1204),
    .Y(_00304_));
 inv_2 _23170_ (.A(net1210),
    .Y(_00305_));
 inv_2 _23171_ (.A(net1208),
    .Y(_00306_));
 inv_2 _23172_ (.A(net1208),
    .Y(_00307_));
 inv_2 _23173_ (.A(net1209),
    .Y(_00308_));
 inv_2 _23174_ (.A(net1206),
    .Y(_00309_));
 inv_2 _23175_ (.A(net1202),
    .Y(_00310_));
 inv_2 _23176_ (.A(net1210),
    .Y(_00311_));
 inv_2 _23177_ (.A(net1202),
    .Y(_00312_));
 inv_2 _23178_ (.A(net1202),
    .Y(_00313_));
 inv_2 _23179_ (.A(net1210),
    .Y(_00314_));
 inv_2 _23180_ (.A(net1207),
    .Y(_00315_));
 inv_2 _23181_ (.A(net1206),
    .Y(_00316_));
 inv_2 _23182_ (.A(net1210),
    .Y(_00317_));
 inv_2 _23183_ (.A(net1201),
    .Y(_00318_));
 inv_2 _23184_ (.A(net1213),
    .Y(_00319_));
 inv_2 _23185_ (.A(net1204),
    .Y(_00320_));
 inv_2 _23186_ (.A(net1213),
    .Y(_00321_));
 inv_2 _23187_ (.A(net1201),
    .Y(_00322_));
 inv_2 _23188_ (.A(net1202),
    .Y(_00323_));
 inv_2 _23189_ (.A(net1213),
    .Y(_00324_));
 inv_2 _23190_ (.A(net1213),
    .Y(_00325_));
 inv_2 _23191_ (.A(net1213),
    .Y(_00326_));
 inv_2 _23192_ (.A(net1213),
    .Y(_00327_));
 inv_2 _23193_ (.A(net1697),
    .Y(_00328_));
 inv_2 _23194_ (.A(net1697),
    .Y(_00329_));
 inv_2 _23195_ (.A(net1202),
    .Y(_00330_));
 inv_2 _23196_ (.A(net1201),
    .Y(_00331_));
 inv_2 _23197_ (.A(net1201),
    .Y(_00332_));
 inv_2 _23198_ (.A(net1202),
    .Y(_00333_));
 inv_2 _23199_ (.A(net1201),
    .Y(_00334_));
 inv_2 _23200_ (.A(net1209),
    .Y(_00335_));
 inv_2 _23201_ (.A(net1205),
    .Y(_00336_));
 inv_2 _23202_ (.A(net1209),
    .Y(_00337_));
 inv_2 _23203_ (.A(net1209),
    .Y(_00338_));
 inv_2 _23204_ (.A(net1209),
    .Y(_00339_));
 inv_2 _23205_ (.A(net1209),
    .Y(_00340_));
 inv_2 _23206_ (.A(net1209),
    .Y(_00341_));
 inv_2 _23207_ (.A(net1211),
    .Y(_00342_));
 inv_2 _23208_ (.A(net1212),
    .Y(_00343_));
 inv_2 _23209_ (.A(net1209),
    .Y(_00344_));
 inv_2 _23210_ (.A(net1209),
    .Y(_00345_));
 inv_2 _23211_ (.A(net1210),
    .Y(_00346_));
 inv_2 _23212_ (.A(net1211),
    .Y(_00347_));
 inv_2 _23213_ (.A(net1210),
    .Y(_00348_));
 or4_1 _23214_ (.A(net1678),
    .B(net1277),
    .C(net1669),
    .D(net1675),
    .X(_00349_));
 or4_1 _23215_ (.A(net1678),
    .B(net1277),
    .C(net1669),
    .D(net1675),
    .X(_00350_));
 or4_1 _23216_ (.A(net1678),
    .B(net1277),
    .C(net1669),
    .D(net1675),
    .X(_00351_));
 or4_1 _23217_ (.A(net1678),
    .B(net1277),
    .C(net1279),
    .D(net1675),
    .X(_00352_));
 dfrtp_1 _23218_ (.CLK(tclk_i),
    .D(_00353_),
    .RESET_B(net1402),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.reg_wr_en ));
 dfrtp_1 _23219_ (.CLK(clk_i),
    .D(ff_erase_after_buf),
    .RESET_B(net1508),
    .Q(ff_erase_ff));
 dfrtp_1 _23220_ (.CLK(clk_i),
    .D(net1815),
    .RESET_B(net1508),
    .Q(ff_erase_ff2));
 dfrtp_1 _23221_ (.CLK(clk_i),
    .D(net1823),
    .RESET_B(net1508),
    .Q(ff_erase_ff3));
 dfrtp_1 _23222_ (.CLK(clk_i),
    .D(ff_prog_after_buf),
    .RESET_B(net1505),
    .Q(ff_prog_ff));
 dfrtp_1 _23223_ (.CLK(clk_i),
    .D(net1810),
    .RESET_B(net1505),
    .Q(ff_prog_ff2));
 dfrtp_1 _23224_ (.CLK(clk_i),
    .D(net1822),
    .RESET_B(net1505),
    .Q(ff_prog_ff3));
 dfrtp_1 _23225_ (.CLK(clk_i),
    .D(net1836),
    .RESET_B(net1579),
    .Q(\digitop_pav2.sl_i ));
 dfrtp_1 _23226_ (.CLK(clk_i),
    .D(net1831),
    .RESET_B(net1579),
    .Q(\digitop_pav2.s3_i ));
 dfrtp_1 _23227_ (.CLK(clk_i),
    .D(net1834),
    .RESET_B(net1581),
    .Q(\digitop_pav2.s2_i ));
 dfrtp_1 _23228_ (.CLK(clk_i),
    .D(s1_set_after_buf),
    .RESET_B(net1579),
    .Q(s1_set_ff));
 dfrtp_1 _23229_ (.CLK(clk_i),
    .D(net1819),
    .RESET_B(net1579),
    .Q(s1_set_ff2));
 dfrtp_1 _23230_ (.CLK(clk_i),
    .D(s1_rst_after_buf),
    .RESET_B(net1579),
    .Q(s1_rst_ff));
 dfrtp_1 _23231_ (.CLK(clk_i),
    .D(net1820),
    .RESET_B(net1580),
    .Q(s1_rst_ff2));
 dfrtp_1 _23232_ (.CLK(clk_i),
    .D(s2_set_after_buf),
    .RESET_B(net1580),
    .Q(s2_set_ff));
 dfrtp_1 _23233_ (.CLK(clk_i),
    .D(net1818),
    .RESET_B(net1580),
    .Q(s2_set_ff2));
 dfrtp_1 _23234_ (.CLK(clk_i),
    .D(s2_rst_after_buf),
    .RESET_B(net1580),
    .Q(s2_rst_ff));
 dfrtp_1 _23235_ (.CLK(clk_i),
    .D(net1811),
    .RESET_B(net1580),
    .Q(s2_rst_ff2));
 dfrtp_1 _23236_ (.CLK(clk_i),
    .D(s3_set_after_buf),
    .RESET_B(net1580),
    .Q(s3_set_ff));
 dfrtp_1 _23237_ (.CLK(clk_i),
    .D(net1813),
    .RESET_B(net1580),
    .Q(s3_set_ff2));
 dfrtp_1 _23238_ (.CLK(clk_i),
    .D(s3_rst_after_buf),
    .RESET_B(net1579),
    .Q(s3_rst_ff));
 dfrtp_1 _23239_ (.CLK(clk_i),
    .D(net1812),
    .RESET_B(net1580),
    .Q(s3_rst_ff2));
 dfrtp_1 _23240_ (.CLK(clk_i),
    .D(sl_set_after_buf),
    .RESET_B(net1579),
    .Q(sl_set_ff));
 dfrtp_1 _23241_ (.CLK(clk_i),
    .D(net1821),
    .RESET_B(net1579),
    .Q(sl_set_ff2));
 dfrtp_1 _23242_ (.CLK(clk_i),
    .D(sl_rst_after_buf),
    .RESET_B(net1579),
    .Q(sl_rst_ff));
 dfrtp_1 _23243_ (.CLK(clk_i),
    .D(net1814),
    .RESET_B(net1579),
    .Q(sl_rst_ff2));
 dfstp_1 _23244_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_00006_),
    .SET_B(net1267),
    .Q(\digitop_pav2.ack_inst.state_ff[0] ));
 dfrtp_1 _23245_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_00040_),
    .RESET_B(net1264),
    .Q(\digitop_pav2.ack_inst.state_ff[1] ));
 dfrtp_1 _23246_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_00041_),
    .RESET_B(net1267),
    .Q(\digitop_pav2.ack_inst.state_ff[2] ));
 dfrtp_2 _23247_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_00042_),
    .RESET_B(net1264),
    .Q(\digitop_pav2.ack_inst.nvm_ack_rd_stb_o ));
 dfxtp_1 _23248_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00000_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[0] ));
 dfxtp_1 _23249_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00001_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[1] ));
 dfxtp_1 _23250_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00002_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[2] ));
 dfxtp_1 _23251_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00003_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[3] ));
 dfxtp_1 _23252_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00004_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[4] ));
 dfxtp_1 _23253_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00005_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[5] ));
 dfstp_1 _23254_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00043_),
    .SET_B(net1437),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[0] ));
 dfrtp_1 _23255_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00044_),
    .RESET_B(net1437),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[1] ));
 dfrtp_2 _23256_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00045_),
    .RESET_B(net1437),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[2] ));
 dfrtp_1 _23257_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00046_),
    .RESET_B(net1437),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[3] ));
 dfrtp_4 _23258_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00047_),
    .RESET_B(net1437),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[4] ));
 dfrtp_4 _23259_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00048_),
    .RESET_B(net1437),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[5] ));
 dfrtp_1 _23260_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00049_),
    .RESET_B(net1444),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[6] ));
 dfrtp_1 _23261_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00050_),
    .RESET_B(net1437),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[7] ));
 dfxtp_4 _23262_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00357_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[0] ));
 dfxtp_4 _23263_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00358_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[1] ));
 dfxtp_2 _23264_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00359_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[2] ));
 dfxtp_2 _23265_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00360_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[3] ));
 dfxtp_2 _23266_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00361_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[4] ));
 dfxtp_2 _23267_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00362_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[5] ));
 dfxtp_2 _23268_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00363_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[6] ));
 dfxtp_4 _23269_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00364_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[7] ));
 dfrtp_1 _23270_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00365_),
    .RESET_B(_00171_),
    .Q(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[6] ));
 dfrtp_1 _23271_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00366_),
    .RESET_B(_00172_),
    .Q(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[4] ));
 dfrtp_1 _23272_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00367_),
    .RESET_B(_00173_),
    .Q(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[5] ));
 dfrtp_1 _23273_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00368_),
    .RESET_B(_00174_),
    .Q(\digitop_pav2.access_inst.access_proc0.proc_crc_check[2] ));
 dfrtp_1 _23274_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00369_),
    .RESET_B(_00175_),
    .Q(\digitop_pav2.access_inst.access_proc0.proc_crc_check[3] ));
 dfrtp_1 _23275_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00370_),
    .RESET_B(_00176_),
    .Q(\digitop_pav2.access_inst.access_proc0.proc_crc_check[4] ));
 dfxtp_1 _23276_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00371_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[1] ));
 dfxtp_1 _23277_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00372_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[2] ));
 dfxtp_1 _23278_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00373_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[3] ));
 dfxtp_1 _23279_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00374_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[4] ));
 dfxtp_1 _23280_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00375_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[5] ));
 dfxtp_1 _23281_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00376_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[6] ));
 dfxtp_1 _23282_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00377_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[7] ));
 dfxtp_1 _23283_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00378_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[8] ));
 dfxtp_1 _23284_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00379_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[9] ));
 dfxtp_1 _23285_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00380_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[10] ));
 dfxtp_1 _23286_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00381_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[11] ));
 dfxtp_1 _23287_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00382_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[12] ));
 dfxtp_1 _23288_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00383_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[13] ));
 dfxtp_1 _23289_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00384_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[14] ));
 dfxtp_1 _23290_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00385_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[15] ));
 dfxtp_1 _23291_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00386_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.txrx_dt_buf[0] ));
 dfxtp_2 _23292_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00387_),
    .Q(\digitop_pav2.access_inst.access_check0.wordcnt_i[0] ));
 dfxtp_2 _23293_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00388_),
    .Q(\digitop_pav2.access_inst.access_check0.wordcnt_i[1] ));
 dfxtp_1 _23294_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00389_),
    .Q(\digitop_pav2.access_inst.access_check0.wordcnt_i[2] ));
 dfxtp_2 _23295_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00390_),
    .Q(\digitop_pav2.access_inst.access_check0.wordcnt_i[3] ));
 dfxtp_1 _23296_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00391_),
    .Q(\digitop_pav2.access_inst.access_check0.wordcnt_i[4] ));
 dfxtp_1 _23297_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00392_),
    .Q(\digitop_pav2.access_inst.access_check0.wordcnt_i[5] ));
 dfxtp_1 _23298_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00393_),
    .Q(\digitop_pav2.access_inst.access_check0.wordcnt_i[6] ));
 dfxtp_1 _23299_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00394_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.rx_par_buf[14] ));
 dfxtp_1 _23300_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00395_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.rx_par_buf[15] ));
 dfxtp_4 _23301_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00396_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[0] ));
 dfxtp_4 _23302_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00397_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[1] ));
 dfxtp_4 _23303_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00398_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[2] ));
 dfxtp_2 _23304_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00399_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[3] ));
 dfxtp_2 _23305_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00400_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[4] ));
 dfxtp_4 _23306_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00401_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[5] ));
 dfxtp_4 _23307_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00402_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[6] ));
 dfxtp_4 _23308_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00403_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[7] ));
 dfxtp_4 _23309_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00404_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[8] ));
 dfxtp_2 _23310_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00405_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[9] ));
 dfxtp_4 _23311_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00406_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ));
 dfxtp_2 _23312_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00407_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[11] ));
 dfxtp_2 _23313_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00408_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[12] ));
 dfxtp_2 _23314_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00409_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[13] ));
 dfxtp_4 _23315_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00410_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[14] ));
 dfxtp_4 _23316_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00411_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[15] ));
 dfxtp_2 _23317_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00412_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[8] ));
 dfxtp_2 _23318_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00413_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[9] ));
 dfxtp_4 _23319_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00414_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[10] ));
 dfxtp_2 _23320_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00415_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[11] ));
 dfxtp_2 _23321_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00416_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[12] ));
 dfxtp_2 _23322_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00417_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[13] ));
 dfxtp_2 _23323_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00418_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[14] ));
 dfxtp_2 _23324_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00419_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[15] ));
 dfxtp_4 _23325_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00420_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[8] ));
 dfxtp_4 _23326_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00421_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[9] ));
 dfxtp_4 _23327_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00422_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ));
 dfxtp_2 _23328_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00423_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[11] ));
 dfxtp_4 _23329_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00424_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[12] ));
 dfxtp_2 _23330_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00425_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[13] ));
 dfxtp_4 _23331_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00426_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[14] ));
 dfxtp_4 _23332_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00427_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[15] ));
 dfxtp_4 _23333_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00428_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[0] ));
 dfxtp_4 _23334_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00429_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[1] ));
 dfxtp_2 _23335_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00430_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[2] ));
 dfxtp_2 _23336_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00431_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[3] ));
 dfxtp_2 _23337_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00432_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[4] ));
 dfxtp_2 _23338_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00433_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[5] ));
 dfxtp_2 _23339_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00434_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[6] ));
 dfxtp_4 _23340_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00435_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[7] ));
 dfxtp_2 _23341_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00436_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[0] ));
 dfxtp_2 _23342_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00437_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[1] ));
 dfxtp_4 _23343_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00438_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[2] ));
 dfxtp_2 _23344_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00439_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[3] ));
 dfxtp_2 _23345_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00440_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[4] ));
 dfxtp_2 _23346_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00441_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[5] ));
 dfxtp_4 _23347_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00442_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[6] ));
 dfxtp_4 _23348_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00443_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ));
 dfxtp_2 _23349_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00444_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[8] ));
 dfxtp_2 _23350_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00445_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[9] ));
 dfxtp_2 _23351_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00446_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[10] ));
 dfxtp_2 _23352_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00447_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[11] ));
 dfxtp_4 _23353_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00448_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[12] ));
 dfxtp_2 _23354_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00449_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[13] ));
 dfxtp_2 _23355_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00450_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[14] ));
 dfxtp_4 _23356_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00451_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[15] ));
 dfrtp_1 _23357_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00452_),
    .RESET_B(net1431),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[0] ));
 dfrtp_1 _23358_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00453_),
    .RESET_B(net1446),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[1] ));
 dfrtp_1 _23359_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00454_),
    .RESET_B(net1432),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[2] ));
 dfrtp_2 _23360_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00455_),
    .RESET_B(net1431),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[3] ));
 dfrtp_1 _23361_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00456_),
    .RESET_B(net1446),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[4] ));
 dfrtp_1 _23362_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00457_),
    .RESET_B(net1432),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[5] ));
 dfrtp_1 _23363_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00458_),
    .RESET_B(net1434),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[6] ));
 dfrtp_1 _23364_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00459_),
    .RESET_B(net1445),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[7] ));
 dfrtp_1 _23365_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00460_),
    .RESET_B(net1436),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[8] ));
 dfrtp_1 _23366_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00461_),
    .RESET_B(net1445),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[9] ));
 dfrtp_1 _23367_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00462_),
    .RESET_B(net1434),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[10] ));
 dfrtp_1 _23368_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00463_),
    .RESET_B(net1434),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[11] ));
 dfstp_1 _23369_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00464_),
    .SET_B(net1435),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[12] ));
 dfrtp_1 _23370_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00465_),
    .RESET_B(net1446),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[13] ));
 dfrtp_1 _23371_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00466_),
    .RESET_B(net1434),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[14] ));
 dfstp_1 _23372_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00467_),
    .SET_B(net1445),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[15] ));
 dfxtp_2 _23373_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00468_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[6] ));
 dfxtp_2 _23374_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00469_),
    .Q(\digitop_pav2.dr ));
 dfxtp_1 _23375_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00470_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[1] ));
 dfxtp_1 _23376_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00471_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[2] ));
 dfxtp_2 _23377_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00472_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[3] ));
 dfxtp_1 _23378_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00473_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[4] ));
 dfxtp_1 _23379_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00474_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[5] ));
 dfxtp_1 _23380_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00475_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[1] ));
 dfxtp_1 _23381_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00476_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[7] ));
 dfxtp_1 _23382_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00477_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[6] ));
 dfxtp_1 _23383_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00478_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[5] ));
 dfxtp_1 _23384_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00479_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[4] ));
 dfxtp_1 _23385_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00480_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[3] ));
 dfxtp_1 _23386_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00481_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[2] ));
 dfxtp_1 _23387_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00482_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[6] ));
 dfxtp_1 _23388_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00483_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[0] ));
 dfxtp_1 _23389_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00484_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[1] ));
 dfxtp_1 _23390_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00485_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[2] ));
 dfxtp_1 _23391_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00486_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[3] ));
 dfxtp_1 _23392_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00487_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[4] ));
 dfxtp_1 _23393_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00488_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[5] ));
 dfrtp_1 _23394_ (.CLK(clk_i),
    .D(net1838),
    .RESET_B(net1580),
    .Q(\digitop_pav2.s1_i ));
 dfstp_1 _23395_ (.CLK(tclk_i),
    .D(_00012_),
    .SET_B(net1410),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[0] ));
 dfrtp_1 _23396_ (.CLK(tclk_i),
    .D(_00116_),
    .RESET_B(net1410),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[1] ));
 dfrtp_1 _23397_ (.CLK(tclk_i),
    .D(_00117_),
    .RESET_B(net1409),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[2] ));
 dfrtp_1 _23398_ (.CLK(tclk_i),
    .D(_00118_),
    .RESET_B(net1409),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[3] ));
 dfrtp_1 _23399_ (.CLK(tclk_i),
    .D(_00119_),
    .RESET_B(net1410),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[4] ));
 dfrtp_1 _23400_ (.CLK(tclk_i),
    .D(_00120_),
    .RESET_B(net1410),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[5] ));
 dfrtp_1 _23401_ (.CLK(tclk_i),
    .D(_00121_),
    .RESET_B(net1410),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[6] ));
 dfrtp_1 _23402_ (.CLK(tclk_i),
    .D(_00122_),
    .RESET_B(net1410),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[7] ));
 dfrtp_1 _23403_ (.CLK(tclk_i),
    .D(_00123_),
    .RESET_B(net1410),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.state[8] ));
 dfstp_1 _23404_ (.CLK(tclk_i),
    .D(_00013_),
    .SET_B(net1403),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[0] ));
 dfrtp_1 _23405_ (.CLK(tclk_i),
    .D(_00124_),
    .RESET_B(net1402),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[2] ));
 dfrtp_4 _23406_ (.CLK(tclk_i),
    .D(_00125_),
    .RESET_B(net1412),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[3] ));
 dfstp_1 _23407_ (.CLK(tclk_i),
    .D(_00011_),
    .SET_B(net1406),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[0] ));
 dfrtp_1 _23408_ (.CLK(tclk_i),
    .D(_00104_),
    .RESET_B(net1406),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_form_end ));
 dfrtp_1 _23409_ (.CLK(tclk_i),
    .D(_00105_),
    .RESET_B(net1405),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[2] ));
 dfrtp_1 _23410_ (.CLK(tclk_i),
    .D(_00106_),
    .RESET_B(net1405),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[3] ));
 dfrtp_1 _23411_ (.CLK(tclk_i),
    .D(_00107_),
    .RESET_B(net1405),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[4] ));
 dfrtp_1 _23412_ (.CLK(tclk_i),
    .D(_00108_),
    .RESET_B(net1406),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[5] ));
 dfrtp_1 _23413_ (.CLK(tclk_i),
    .D(_00109_),
    .RESET_B(net1406),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[6] ));
 dfrtp_1 _23414_ (.CLK(tclk_i),
    .D(_00110_),
    .RESET_B(net1406),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[7] ));
 dfrtp_1 _23415_ (.CLK(tclk_i),
    .D(_00111_),
    .RESET_B(net1406),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.state[8] ));
 dfstp_1 _23416_ (.CLK(tclk_i),
    .D(_00112_),
    .SET_B(net1409),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[0] ));
 dfrtp_1 _23417_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_state[2] ),
    .RESET_B(net1415),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[1] ));
 dfrtp_4 _23418_ (.CLK(tclk_i),
    .D(_00113_),
    .RESET_B(net1415),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[2] ));
 dfrtp_1 _23419_ (.CLK(tclk_i),
    .D(_00114_),
    .RESET_B(net1415),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[3] ));
 dfrtp_1 _23420_ (.CLK(tclk_i),
    .D(_00115_),
    .RESET_B(net1415),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.state[4] ));
 dfstp_1 _23421_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00490_),
    .SET_B(net1005),
    .Q(\digitop_pav2.sec_inst.sm.next_st[1] ));
 dfrtp_1 _23422_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00491_),
    .RESET_B(net1005),
    .Q(\digitop_pav2.sec_inst.sm.st[1] ));
 dfrtp_1 _23423_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00492_),
    .RESET_B(net1621),
    .Q(\digitop_pav2.sec_inst.en_ld_r ));
 dfrtp_2 _23424_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00493_),
    .RESET_B(net1621),
    .Q(\digitop_pav2.rng_inst.rng_prngx_pav2.rngx_sec_req_i ));
 dfrtp_1 _23425_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00494_),
    .RESET_B(net1006),
    .Q(\digitop_pav2.sec_inst.en_ld_data ));
 dfrtp_1 _23426_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(net1648),
    .RESET_B(net1006),
    .Q(\digitop_pav2.sec_inst.dg_key.en_i ));
 dfrtp_2 _23427_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00496_),
    .RESET_B(net1006),
    .Q(\digitop_pav2.sec_inst.sm.st[6] ));
 dfrtp_1 _23428_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00497_),
    .RESET_B(net1006),
    .Q(\digitop_pav2.sec_inst.en_shifto ));
 dfrtp_1 _23429_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00498_),
    .RESET_B(net1006),
    .Q(\digitop_pav2.sec_inst.en_reg128 ));
 dfrtp_4 _23430_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00499_),
    .RESET_B(net1621),
    .Q(\digitop_pav2.sec_inst.sm.st[9] ));
 dfstp_1 _23431_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00008_),
    .SET_B(net986),
    .Q(\digitop_pav2.sec_inst.shift_out.st[0] ));
 dfrtp_1 _23432_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00009_),
    .RESET_B(net986),
    .Q(\digitop_pav2.sec_inst.shift_out.st[2] ));
 dfrtp_1 _23433_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00100_),
    .RESET_B(net984),
    .Q(\digitop_pav2.sec_inst.shift_out.st[3] ));
 dfrtp_1 _23434_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00010_),
    .RESET_B(net985),
    .Q(\digitop_pav2.sec_inst.shift_out.st[4] ));
 dfrtp_1 _23435_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00101_),
    .RESET_B(net986),
    .Q(\digitop_pav2.sec_inst.shift_out.st[5] ));
 dfrtp_1 _23436_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00102_),
    .RESET_B(net985),
    .Q(\digitop_pav2.sec_inst.shift_out.st[6] ));
 dfrtp_1 _23437_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00103_),
    .RESET_B(net986),
    .Q(\digitop_pav2.sec_inst.shift_out.st[7] ));
 dfstp_2 _23438_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00098_),
    .SET_B(net1005),
    .Q(\digitop_pav2.sec_inst.ld_mem.st[0] ));
 dfrtp_1 _23439_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00099_),
    .RESET_B(net1005),
    .Q(\digitop_pav2.sec_inst.ld_mem.st[1] ));
 dfstp_1 _23440_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00082_),
    .SET_B(net1447),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[0] ));
 dfrtp_2 _23441_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00087_),
    .RESET_B(net1449),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[1] ));
 dfrtp_1 _23442_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00088_),
    .RESET_B(net1447),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[2] ));
 dfrtp_1 _23443_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00089_),
    .RESET_B(net1448),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[3] ));
 dfrtp_1 _23444_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00090_),
    .RESET_B(net1448),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[4] ));
 dfrtp_4 _23445_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00091_),
    .RESET_B(net1448),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[5] ));
 dfrtp_1 _23446_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00092_),
    .RESET_B(net1449),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[6] ));
 dfrtp_2 _23447_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00093_),
    .RESET_B(net1448),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[7] ));
 dfrtp_1 _23448_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00094_),
    .RESET_B(net1449),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[8] ));
 dfrtp_1 _23449_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00095_),
    .RESET_B(net1448),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[9] ));
 dfrtp_1 _23450_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00083_),
    .RESET_B(net1448),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.cg_en_13 ));
 dfrtp_2 _23451_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00084_),
    .RESET_B(net1448),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[11] ));
 dfrtp_2 _23452_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00085_),
    .RESET_B(net1448),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[12] ));
 dfrtp_1 _23453_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00086_),
    .RESET_B(net1449),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[13] ));
 dfstp_1 _23454_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_00078_),
    .SET_B(net1420),
    .Q(\digitop_pav2.memctrl_inst.state[0] ));
 dfrtp_1 _23455_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(\digitop_pav2.memctrl_inst.n_state[2] ),
    .RESET_B(net1425),
    .Q(\digitop_pav2.memctrl_inst.state[1] ));
 dfrtp_1 _23456_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_00079_),
    .RESET_B(net1425),
    .Q(\digitop_pav2.memctrl_inst.state[2] ));
 dfrtp_1 _23457_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_00080_),
    .RESET_B(net1419),
    .Q(\digitop_pav2.memctrl_inst.state[3] ));
 dfrtp_1 _23458_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_00081_),
    .RESET_B(net1419),
    .Q(\digitop_pav2.memctrl_inst.state[4] ));
 dfstp_1 _23459_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00014_),
    .SET_B(_00177_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[0] ));
 dfrtp_1 _23460_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00025_),
    .RESET_B(_00178_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[1] ));
 dfrtp_1 _23461_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00032_),
    .RESET_B(_00179_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[2] ));
 dfrtp_1 _23462_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00033_),
    .RESET_B(_00180_),
    .Q(\digitop_pav2.access_inst.access_check0.write_check_i ));
 dfrtp_1 _23463_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00034_),
    .RESET_B(_00181_),
    .Q(\digitop_pav2.access_inst.access_check0.wr_key_ck_i ));
 dfrtp_1 _23464_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00035_),
    .RESET_B(_00182_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[5] ));
 dfrtp_2 _23465_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00036_),
    .RESET_B(_00183_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.crc_en_o ));
 dfrtp_2 _23466_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00037_),
    .RESET_B(_00184_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt_ok ));
 dfrtp_1 _23467_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00038_),
    .RESET_B(_00185_),
    .Q(\digitop_pav2.access_inst.access_check0.pc_lock_check_i ));
 dfrtp_1 _23468_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00039_),
    .RESET_B(_00186_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[9] ));
 dfrtp_1 _23469_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00015_),
    .RESET_B(_00187_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[10] ));
 dfrtp_1 _23470_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00016_),
    .RESET_B(_00188_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[11] ));
 dfrtp_1 _23471_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00017_),
    .RESET_B(_00189_),
    .Q(\digitop_pav2.access_inst.access_check0.mem_sign_check_i ));
 dfrtp_2 _23472_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00018_),
    .RESET_B(_00190_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[13] ));
 dfrtp_1 _23473_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00019_),
    .RESET_B(_00191_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[14] ));
 dfrtp_1 _23474_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00020_),
    .RESET_B(_00192_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[15] ));
 dfrtp_2 _23475_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00021_),
    .RESET_B(_00193_),
    .Q(\digitop_pav2.access_inst.access_check0.wr_lock_ck_i ));
 dfrtp_1 _23476_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00022_),
    .RESET_B(_00194_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[17] ));
 dfrtp_1 _23477_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00023_),
    .RESET_B(_00195_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[18] ));
 dfrtp_1 _23478_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00024_),
    .RESET_B(_00196_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[19] ));
 dfrtp_1 _23479_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00026_),
    .RESET_B(_00197_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[20] ));
 dfrtp_4 _23480_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00027_),
    .RESET_B(_00198_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.ld_dt_stb ));
 dfrtp_1 _23481_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00028_),
    .RESET_B(_00199_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[22] ));
 dfrtp_1 _23482_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00029_),
    .RESET_B(_00200_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[23] ));
 dfrtp_1 _23483_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00030_),
    .RESET_B(_00201_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[24] ));
 dfrtp_1 _23484_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_00031_),
    .RESET_B(_00202_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.state[25] ));
 dfrtp_1 _23485_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00096_),
    .RESET_B(net972),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[4] ));
 dfrtp_1 _23486_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00097_),
    .RESET_B(net972),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[8] ));
 dfrtp_1 _23487_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_state[0] ),
    .RESET_B(net1403),
    .Q(\digitop_pav2.testctrl_pav2.inst_mode.state[0] ));
 dfrtp_1 _23488_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_state[1] ),
    .RESET_B(net1404),
    .Q(\digitop_pav2.testctrl_pav2.inst_mode.state[1] ));
 dfrtp_1 _23489_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_state[2] ),
    .RESET_B(net1403),
    .Q(\digitop_pav2.testctrl_pav2.inst_mode.state[2] ));
 dfrtp_1 _23490_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_state[3] ),
    .RESET_B(net1403),
    .Q(\digitop_pav2.testctrl_pav2.inst_mode.state[3] ));
 dfrtp_1 _23491_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_state[4] ),
    .RESET_B(net1404),
    .Q(\digitop_pav2.testctrl_pav2.inst_mode.state[4] ));
 dfrtp_1 _23492_ (.CLK(\digitop_pav2.sync_inst.inst_rstx.osc_clk_gated ),
    .D(_00500_),
    .RESET_B(\digitop_pav2.sync_inst.inst_rstx.sync_rstx_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.sync_inst.inst_rstx.gray_counter[1] ));
 dfrtp_1 _23493_ (.CLK(\digitop_pav2.sync_inst.inst_rstx.osc_clk_gated ),
    .D(_00501_),
    .RESET_B(\digitop_pav2.sync_inst.inst_rstx.sync_rstx_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.sync_inst.inst_rstx.gray_counter[2] ));
 dfrtp_1 _23494_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_calclk ),
    .RESET_B(net1403),
    .Q(\digitop_pav2.cal_inst.calx_mux.en_calx_test_i ));
 dfrtp_1 _23495_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_digfunc ),
    .RESET_B(net1403),
    .Q(\digitop_pav2.testctrl_pav2.inst_mode.tm_digfunc ));
 dfrtp_1 _23496_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_anafunc ),
    .RESET_B(net1404),
    .Q(\digitop_pav2.testctrl_pav2.inst_mode.tm_anafunc ));
 dfrtp_1 _23497_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_probe ),
    .RESET_B(net1403),
    .Q(\digitop_pav2.testctrl_pav2.inst_mode.tm_probe ));
 dfrtp_1 _23498_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_dummy ),
    .RESET_B(net1403),
    .Q(\digitop_pav2.testctrl_pav2.inst_mode.tm_dummy ));
 dfrtp_1 _23499_ (.CLK(tclk_i),
    .D(_00162_),
    .RESET_B(net1402),
    .Q(\digitop_pav2.testctrl_pav2.inst_mode.tm_amux ));
 dfrtp_4 _23500_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_rnclkout ),
    .RESET_B(net1403),
    .Q(\digitop_pav2.testctrl_pav2.inst_mode.tm_rnclkout ));
 dfrtp_2 _23501_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_clkout ),
    .RESET_B(net1404),
    .Q(\digitop_pav2.testctrl_pav2.inst_mode.tm_clkout ));
 dfrtp_4 _23502_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mode.n_tm_mbist ),
    .RESET_B(net1403),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.tm_mbist_i ));
 dfrtp_1 _23503_ (.CLK(tclk_i),
    .D(_00165_),
    .RESET_B(net1401),
    .Q(\digitop_pav2.testctrl_pav2.inst_tmamux.window_vcc ));
 dfrtp_1 _23504_ (.CLK(tclk_i),
    .D(_00167_),
    .RESET_B(net1402),
    .Q(\digitop_pav2.testctrl_pav2.inst_tmamux.window_vref ));
 dfrtp_1 _23505_ (.CLK(tclk_i),
    .D(_00166_),
    .RESET_B(net1401),
    .Q(\digitop_pav2.testctrl_pav2.inst_tmamux.window_vdd ));
 dfrtp_1 _23506_ (.CLK(tclk_i),
    .D(_00164_),
    .RESET_B(net1401),
    .Q(\digitop_pav2.testctrl_pav2.inst_tmamux.window_ibias ));
 dfrtp_1 _23507_ (.CLK(_00203_),
    .D(_00163_),
    .RESET_B(net1402),
    .Q(net70));
 dfstp_1 _23508_ (.CLK(tclk_i),
    .D(_00502_),
    .SET_B(net1411),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[0] ));
 dfstp_1 _23509_ (.CLK(tclk_i),
    .D(_00503_),
    .SET_B(net1411),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[1] ));
 dfstp_1 _23510_ (.CLK(tclk_i),
    .D(_00504_),
    .SET_B(net1411),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[2] ));
 dfstp_1 _23511_ (.CLK(tclk_i),
    .D(_00505_),
    .SET_B(net1411),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[3] ));
 dfstp_1 _23512_ (.CLK(tclk_i),
    .D(_00506_),
    .SET_B(net1409),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[4] ));
 dfstp_1 _23513_ (.CLK(tclk_i),
    .D(_00507_),
    .SET_B(net1411),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.ctr[5] ));
 dfrtp_1 _23514_ (.CLK(tclk_i),
    .D(_00508_),
    .RESET_B(net1422),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[0] ));
 dfrtp_1 _23515_ (.CLK(tclk_i),
    .D(_00509_),
    .RESET_B(net1422),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[1] ));
 dfrtp_1 _23516_ (.CLK(tclk_i),
    .D(_00510_),
    .RESET_B(net1422),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[2] ));
 dfrtp_1 _23517_ (.CLK(tclk_i),
    .D(_00511_),
    .RESET_B(net1422),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[3] ));
 dfrtp_1 _23518_ (.CLK(tclk_i),
    .D(_00512_),
    .RESET_B(net1422),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[4] ));
 dfrtp_1 _23519_ (.CLK(tclk_i),
    .D(_00513_),
    .RESET_B(net1422),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[5] ));
 dfrtp_1 _23520_ (.CLK(tclk_i),
    .D(_00514_),
    .RESET_B(net1422),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[6] ));
 dfrtp_1 _23521_ (.CLK(tclk_i),
    .D(_00515_),
    .RESET_B(net1423),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[7] ));
 dfrtp_1 _23522_ (.CLK(tclk_i),
    .D(_00516_),
    .RESET_B(net1423),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[8] ));
 dfrtp_1 _23523_ (.CLK(tclk_i),
    .D(_00517_),
    .RESET_B(net1423),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[9] ));
 dfrtp_1 _23524_ (.CLK(tclk_i),
    .D(_00518_),
    .RESET_B(net1423),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[10] ));
 dfrtp_1 _23525_ (.CLK(tclk_i),
    .D(_00519_),
    .RESET_B(net1423),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[11] ));
 dfrtp_1 _23526_ (.CLK(tclk_i),
    .D(_00520_),
    .RESET_B(net1422),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[12] ));
 dfrtp_1 _23527_ (.CLK(tclk_i),
    .D(_00521_),
    .RESET_B(net1422),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[13] ));
 dfrtp_1 _23528_ (.CLK(tclk_i),
    .D(_00522_),
    .RESET_B(net1423),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[14] ));
 dfrtp_2 _23529_ (.CLK(tclk_i),
    .D(_00523_),
    .RESET_B(net1423),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[15] ));
 dfrtp_1 _23530_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_prog ),
    .RESET_B(net1416),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.rr_prog ));
 dfstp_1 _23531_ (.CLK(tclk_i),
    .D(_00524_),
    .SET_B(net1405),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[0] ));
 dfstp_1 _23532_ (.CLK(tclk_i),
    .D(_00525_),
    .SET_B(net1405),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[1] ));
 dfstp_1 _23533_ (.CLK(tclk_i),
    .D(_00526_),
    .SET_B(net1405),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[2] ));
 dfstp_1 _23534_ (.CLK(tclk_i),
    .D(_00527_),
    .SET_B(net1421),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[3] ));
 dfstp_1 _23535_ (.CLK(tclk_i),
    .D(_00528_),
    .SET_B(net1408),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.wlnum[4] ));
 dfstp_1 _23536_ (.CLK(tclk_i),
    .D(_00529_),
    .SET_B(net1416),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[0] ));
 dfstp_1 _23537_ (.CLK(tclk_i),
    .D(_00530_),
    .SET_B(net1416),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[1] ));
 dfstp_1 _23538_ (.CLK(tclk_i),
    .D(_00531_),
    .SET_B(net1419),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[2] ));
 dfstp_1 _23539_ (.CLK(tclk_i),
    .D(_00532_),
    .SET_B(net1421),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.bitctr[3] ));
 dfrtp_4 _23540_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_int_wr_end ),
    .RESET_B(net1409),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_end_i ));
 dfrtp_1 _23541_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_read ),
    .RESET_B(net1415),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.rr_read ));
 dfrtp_1 _23542_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_int_rd_end ),
    .RESET_B(net1411),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rd_end_i ));
 dfrtp_1 _23543_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.n_rr_erase ),
    .RESET_B(net1416),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.rr_erase ));
 dfrtp_1 _23544_ (.CLK(tclk_i),
    .D(_00533_),
    .RESET_B(net1414),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[0] ));
 dfrtp_1 _23545_ (.CLK(tclk_i),
    .D(_00534_),
    .RESET_B(net1421),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[1] ));
 dfrtp_1 _23546_ (.CLK(tclk_i),
    .D(_00535_),
    .RESET_B(net1414),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[2] ));
 dfrtp_1 _23547_ (.CLK(tclk_i),
    .D(_00536_),
    .RESET_B(net1414),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[3] ));
 dfrtp_2 _23548_ (.CLK(tclk_i),
    .D(_00537_),
    .RESET_B(net1414),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[4] ));
 dfrtp_1 _23549_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.n_int_wr_stb ),
    .RESET_B(net1405),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.int_wr_stb ));
 dfrtp_1 _23550_ (.CLK(tclk_i),
    .D(_00538_),
    .RESET_B(net1410),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.mbist_end ));
 dfrtp_2 _23551_ (.CLK(tclk_i),
    .D(_00539_),
    .RESET_B(net1410),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.mbist_result ));
 dfrtp_1 _23552_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.n_int_wr_bit ),
    .RESET_B(net1405),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.int_wr_bit ));
 dfrtp_1 _23553_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.n_int_rd_stb ),
    .RESET_B(net1409),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.int_rd_stb ));
 dfrtp_1 _23554_ (.CLK(tclk_i),
    .D(_00540_),
    .RESET_B(net1406),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.read_after_prog_ok ));
 dfrtp_1 _23555_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_form_enable ),
    .RESET_B(net1406),
    .Q(net105));
 dfrtp_1 _23556_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_int_wr_stb ),
    .RESET_B(net1405),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_stb ));
 dfstp_1 _23557_ (.CLK(tclk_i),
    .D(_00541_),
    .SET_B(net1407),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[0] ));
 dfstp_1 _23558_ (.CLK(tclk_i),
    .D(_00542_),
    .SET_B(net1407),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[1] ));
 dfstp_1 _23559_ (.CLK(tclk_i),
    .D(_00543_),
    .SET_B(net1407),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[2] ));
 dfstp_1 _23560_ (.CLK(tclk_i),
    .D(_00544_),
    .SET_B(net1407),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[3] ));
 dfstp_1 _23561_ (.CLK(tclk_i),
    .D(_00545_),
    .SET_B(net1407),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[4] ));
 dfstp_1 _23562_ (.CLK(tclk_i),
    .D(_00546_),
    .SET_B(net1407),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[5] ));
 dfstp_1 _23563_ (.CLK(tclk_i),
    .D(_00547_),
    .SET_B(net1407),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[6] ));
 dfstp_1 _23564_ (.CLK(tclk_i),
    .D(_00548_),
    .SET_B(net1407),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[7] ));
 dfstp_1 _23565_ (.CLK(tclk_i),
    .D(_00549_),
    .SET_B(net1407),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[8] ));
 dfstp_1 _23566_ (.CLK(tclk_i),
    .D(_00550_),
    .SET_B(net1406),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.ctr[9] ));
 dfrtp_1 _23567_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_form_end ),
    .RESET_B(net1406),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.form_end ));
 dfrtp_1 _23568_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_int_wr_bit ),
    .RESET_B(net1408),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_wr_bit ));
 dfrtp_1 _23569_ (.CLK(tclk_i),
    .D(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.n_int_rd_stb ),
    .RESET_B(net1409),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rd_stb ));
 dfrtp_1 _23570_ (.CLK(\digitop_pav2.testctrl_pav2.inst_enter.tmrboot_clk ),
    .D(_00551_),
    .RESET_B(net1404),
    .Q(\digitop_pav2.testctrl_pav2.inst_enter.tm_enter ));
 dfstp_1 _23571_ (.CLK(tclk_i),
    .D(_00552_),
    .SET_B(net1401),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[0] ));
 dfstp_1 _23572_ (.CLK(tclk_i),
    .D(_00553_),
    .SET_B(net1401),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[1] ));
 dfstp_1 _23573_ (.CLK(tclk_i),
    .D(_00554_),
    .SET_B(net1401),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[2] ));
 dfstp_1 _23574_ (.CLK(tclk_i),
    .D(_00555_),
    .SET_B(net1401),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[3] ));
 dfstp_1 _23575_ (.CLK(tclk_i),
    .D(_00556_),
    .SET_B(net1401),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[4] ));
 dfstp_1 _23576_ (.CLK(tclk_i),
    .D(_00557_),
    .SET_B(net1401),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[5] ));
 dfstp_1 _23577_ (.CLK(tclk_i),
    .D(_00558_),
    .SET_B(net1401),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[6] ));
 dfstp_1 _23578_ (.CLK(tclk_i),
    .D(_00559_),
    .SET_B(net1402),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[7] ));
 dfstp_1 _23579_ (.CLK(tclk_i),
    .D(_00560_),
    .SET_B(net1402),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[8] ));
 dfstp_1 _23580_ (.CLK(tclk_i),
    .D(_00561_),
    .SET_B(net1402),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_regwen.regwctr[9] ));
 dfstp_1 _23581_ (.CLK(tclk_i),
    .D(_00562_),
    .SET_B(net1409),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[0] ));
 dfstp_1 _23582_ (.CLK(tclk_i),
    .D(_00563_),
    .SET_B(net1405),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[1] ));
 dfstp_1 _23583_ (.CLK(tclk_i),
    .D(_00564_),
    .SET_B(net1408),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[2] ));
 dfstp_1 _23584_ (.CLK(tclk_i),
    .D(_00565_),
    .SET_B(net1409),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[3] ));
 dfstp_1 _23585_ (.CLK(tclk_i),
    .D(_00566_),
    .SET_B(net1409),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_mbist.wlnum[4] ));
 dfrtp_1 _23586_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.rngx_pup_clk_i ),
    .D(_00567_),
    .RESET_B(net1442),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[0] ));
 dfrtp_1 _23587_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.rngx_pup_clk_i ),
    .D(_00568_),
    .RESET_B(net1442),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[1] ));
 dfrtp_1 _23588_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.rngx_pup_clk_i ),
    .D(_00569_),
    .RESET_B(net1442),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[2] ));
 dfrtp_1 _23589_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.rngx_pup_clk_i ),
    .D(_00570_),
    .RESET_B(net1442),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[3] ));
 dfrtp_1 _23590_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.rngx_pup_clk_i ),
    .D(_00571_),
    .RESET_B(net1442),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[4] ));
 dfrtp_1 _23591_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.rngx_pup_clk_i ),
    .D(_00572_),
    .RESET_B(net1442),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[5] ));
 dfrtp_1 _23592_ (.CLK(\digitop_pav2.sync_inst.inst_rstx.osc_clk_gated ),
    .D(_00573_),
    .RESET_B(\digitop_pav2.sync_inst.inst_rstx.sync_rstx_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.aes128_inst.aes128_counter.rst_b_i ));
 dfstp_1 _23593_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_fc_clk ),
    .D(_00146_),
    .SET_B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux ),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ));
 dfstp_1 _23594_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.mode_after_buf ),
    .D(net1585),
    .SET_B(_00204_),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.en_blf_fc_b ));
 dfrtp_1 _23595_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk ),
    .D(\digitop_pav2.pass_t2 ),
    .RESET_B(_00205_),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.pass_t2_ff ));
 dfstp_1 _23596_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[5].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .D(_00152_),
    .SET_B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux ),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.A ));
 dfstp_1 _23597_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .D(_00150_),
    .SET_B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux ),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.A ));
 dfstp_1 _23598_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .D(_00153_),
    .SET_B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux ),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[7].sync_pav2_clkx_delay_DONT_TOUCH.A ));
 dfstp_1 _23599_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .D(_00149_),
    .SET_B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux ),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.A ));
 dfstp_1 _23600_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .D(_00148_),
    .SET_B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux ),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.A ));
 dfstp_1 _23601_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .D(_00151_),
    .SET_B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux ),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[5].sync_pav2_clkx_delay_DONT_TOUCH.A ));
 dfstp_1 _23602_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .D(_00147_),
    .SET_B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux ),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.A ));
 dfstp_1 _23603_ (.CLK(_00207_),
    .D(_00155_),
    .SET_B(_00206_),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_mask_before_buf ));
 dfstp_1 _23604_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk ),
    .D(_00574_),
    .SET_B(_00208_),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.dis_blf_fc_b ));
 dfrtp_1 _23605_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_fc_clk_gated ),
    .D(_00154_),
    .RESET_B(_00209_),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.en_ctr ));
 dfstp_1 _23606_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m2_clk_after_buf ),
    .D(_00157_),
    .SET_B(\digitop_pav2.sync_inst.inst_clkx.inst_cp.int_rst_b ),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m4_clk ));
 dfstp_1 _23607_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m4_clk_after_buf ),
    .D(_00158_),
    .SET_B(\digitop_pav2.sync_inst.inst_clkx.inst_cp.int_rst_b ),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m8_clk ));
 dfstp_1 _23608_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.blf_clk ),
    .D(_00575_),
    .SET_B(net1726),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_fm0x.en_fm0x_clk_b ));
 dfstp_1 _23609_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_fc_clk_gated ),
    .D(_00576_),
    .SET_B(_00211_),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk_before_buf ));
 dfstp_1 _23610_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.dft_div4_clk ),
    .D(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_ff.slow_clk_en_b_ff ),
    .SET_B(net1441),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_en.slow_clk_en_b_ff2_i ));
 dfstp_1 _23611_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.dft_div4_clk ),
    .D(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_ff.slow_clk_en_b_i ),
    .SET_B(net1441),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_ff.slow_clk_en_b_ff ));
 dfrtp_1 _23612_ (.CLK(_00212_),
    .D(_00577_),
    .RESET_B(net1436),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_mem.en_mem_clk ));
 dfrtp_1 _23613_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.dft_div4_clk ),
    .D(_00578_),
    .RESET_B(net1441),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div4_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ));
 dfstp_1 _23614_ (.CLK(\digitop_pav2.clkx_piex_clk ),
    .D(\digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_ff2 ),
    .SET_B(net1441),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_ff3 ));
 dfstp_1 _23615_ (.CLK(\digitop_pav2.clkx_piex_clk ),
    .D(\digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_i ),
    .SET_B(net1441),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_ff ));
 dfstp_1 _23616_ (.CLK(\digitop_pav2.clkx_piex_clk ),
    .D(\digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_ff ),
    .SET_B(net1441),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_ff2 ));
 dfstp_1 _23617_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.div2_clk ),
    .D(_00160_),
    .SET_B(net1441),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.div4 ));
 dfstp_1 _23618_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_div4.div_gated_clk ),
    .D(_00159_),
    .SET_B(net1441),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.div2 ));
 dfrtp_1 _23619_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.scwend_clk_i ),
    .D(_00579_),
    .RESET_B(net1442),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.en_scwend_clk_b ));
 dfstp_1 _23620_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.dft_div4_clk ),
    .D(_00580_),
    .SET_B(net1441),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_en.slow_clk_en_b_ff3 ));
 dfstp_1 _23621_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.scwend_clk_i ),
    .D(net1584),
    .SET_B(net1442),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.en_pup_clk_b_aux ));
 dfstp_1 _23622_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.scwend_clk_i ),
    .D(_00581_),
    .SET_B(net1442),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.en_pup_clk_b ));
 dfrtp_1 _23623_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.trigger_clk_i ),
    .D(_00161_),
    .RESET_B(net1442),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.slow_clk_en ));
 dfrtp_1 _23624_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.inst_cgate.ck_in ),
    .D(_00582_),
    .RESET_B(_00213_),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_cipher.inst_en.cipher_off_ff ));
 dfstp_1 _23625_ (.CLK(\digitop_pav2.sync_inst.inst_clkx.blf_clk ),
    .D(_00156_),
    .SET_B(\digitop_pav2.sync_inst.inst_clkx.inst_cp.int_rst_b ),
    .Q(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m2_clk ));
 dfrtp_2 _23626_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00583_),
    .RESET_B(net1005),
    .Q(\digitop_pav2.sec_inst.ld_mem.wctr[0] ));
 dfrtp_2 _23627_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00584_),
    .RESET_B(net1005),
    .Q(\digitop_pav2.sec_inst.ld_mem.wctr[1] ));
 dfrtp_1 _23628_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00585_),
    .RESET_B(net1005),
    .Q(\digitop_pav2.sec_inst.ld_mem.wctr[2] ));
 dfrtp_4 _23629_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00586_),
    .RESET_B(net1005),
    .Q(\digitop_pav2.sec_inst.ld_mem.wctr[3] ));
 dfxtp_2 _23630_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00587_),
    .Q(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[0] ));
 dfxtp_1 _23631_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00588_),
    .Q(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[1] ));
 dfxtp_1 _23632_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00589_),
    .Q(\digitop_pav2.rng_inst.rng_prngx_pav2.sel[2] ));
 dfrtp_4 _23633_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00590_),
    .RESET_B(net1003),
    .Q(\digitop_pav2.sec_inst.ld_r.st[0] ));
 dfrtp_2 _23634_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00591_),
    .RESET_B(net985),
    .Q(\digitop_pav2.sec_inst.ld_r.st[1] ));
 dfstp_1 _23635_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00592_),
    .SET_B(net993),
    .Q(\digitop_pav2.sec_inst.reg160[16] ));
 dfrtp_1 _23636_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00593_),
    .RESET_B(net996),
    .Q(\digitop_pav2.sec_inst.reg160[17] ));
 dfrtp_1 _23637_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00594_),
    .RESET_B(net993),
    .Q(\digitop_pav2.sec_inst.reg160[18] ));
 dfrtp_1 _23638_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00595_),
    .RESET_B(net993),
    .Q(\digitop_pav2.sec_inst.reg160[19] ));
 dfrtp_1 _23639_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00596_),
    .RESET_B(net993),
    .Q(\digitop_pav2.sec_inst.reg160[20] ));
 dfrtp_1 _23640_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00597_),
    .RESET_B(net993),
    .Q(\digitop_pav2.sec_inst.reg160[21] ));
 dfrtp_1 _23641_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00598_),
    .RESET_B(net993),
    .Q(\digitop_pav2.sec_inst.reg160[22] ));
 dfrtp_1 _23642_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00599_),
    .RESET_B(net994),
    .Q(\digitop_pav2.sec_inst.reg160[23] ));
 dfrtp_1 _23643_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00600_),
    .RESET_B(net994),
    .Q(\digitop_pav2.sec_inst.reg160[24] ));
 dfrtp_1 _23644_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00601_),
    .RESET_B(net994),
    .Q(\digitop_pav2.sec_inst.reg160[25] ));
 dfrtp_1 _23645_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00602_),
    .RESET_B(net994),
    .Q(\digitop_pav2.sec_inst.reg160[26] ));
 dfrtp_1 _23646_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00603_),
    .RESET_B(net994),
    .Q(\digitop_pav2.sec_inst.reg160[27] ));
 dfrtp_1 _23647_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00604_),
    .RESET_B(net994),
    .Q(\digitop_pav2.sec_inst.reg160[28] ));
 dfrtp_1 _23648_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00605_),
    .RESET_B(net995),
    .Q(\digitop_pav2.sec_inst.reg160[29] ));
 dfrtp_1 _23649_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00606_),
    .RESET_B(net994),
    .Q(\digitop_pav2.sec_inst.reg160[30] ));
 dfrtp_1 _23650_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00607_),
    .RESET_B(net994),
    .Q(\digitop_pav2.sec_inst.reg160[31] ));
 dfstp_1 _23651_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00608_),
    .SET_B(net996),
    .Q(\digitop_pav2.sec_inst.reg160[32] ));
 dfrtp_1 _23652_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00609_),
    .RESET_B(net995),
    .Q(\digitop_pav2.sec_inst.reg160[33] ));
 dfrtp_1 _23653_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00610_),
    .RESET_B(net995),
    .Q(\digitop_pav2.sec_inst.reg160[34] ));
 dfrtp_1 _23654_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00611_),
    .RESET_B(net995),
    .Q(\digitop_pav2.sec_inst.reg160[35] ));
 dfrtp_1 _23655_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00612_),
    .RESET_B(net995),
    .Q(\digitop_pav2.sec_inst.reg160[36] ));
 dfrtp_1 _23656_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00613_),
    .RESET_B(net994),
    .Q(\digitop_pav2.sec_inst.reg160[37] ));
 dfrtp_1 _23657_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00614_),
    .RESET_B(net998),
    .Q(\digitop_pav2.sec_inst.reg160[38] ));
 dfrtp_1 _23658_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00615_),
    .RESET_B(net998),
    .Q(\digitop_pav2.sec_inst.reg160[39] ));
 dfrtp_1 _23659_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00616_),
    .RESET_B(net998),
    .Q(\digitop_pav2.sec_inst.reg160[40] ));
 dfrtp_1 _23660_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00617_),
    .RESET_B(net998),
    .Q(\digitop_pav2.sec_inst.reg160[41] ));
 dfrtp_1 _23661_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00618_),
    .RESET_B(net998),
    .Q(\digitop_pav2.sec_inst.reg160[42] ));
 dfrtp_1 _23662_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00619_),
    .RESET_B(net998),
    .Q(\digitop_pav2.sec_inst.reg160[43] ));
 dfrtp_1 _23663_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00620_),
    .RESET_B(net998),
    .Q(\digitop_pav2.sec_inst.reg160[44] ));
 dfrtp_1 _23664_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00621_),
    .RESET_B(net997),
    .Q(\digitop_pav2.sec_inst.reg160[45] ));
 dfrtp_1 _23665_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00622_),
    .RESET_B(net997),
    .Q(\digitop_pav2.sec_inst.reg160[46] ));
 dfrtp_1 _23666_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00623_),
    .RESET_B(net997),
    .Q(\digitop_pav2.sec_inst.reg160[47] ));
 dfstp_1 _23667_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00624_),
    .SET_B(net993),
    .Q(\digitop_pav2.sec_inst.reg160[48] ));
 dfrtp_1 _23668_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00625_),
    .RESET_B(net993),
    .Q(\digitop_pav2.sec_inst.reg160[49] ));
 dfrtp_1 _23669_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00626_),
    .RESET_B(net993),
    .Q(\digitop_pav2.sec_inst.reg160[50] ));
 dfrtp_1 _23670_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00627_),
    .RESET_B(net994),
    .Q(\digitop_pav2.sec_inst.reg160[51] ));
 dfrtp_1 _23671_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00628_),
    .RESET_B(net997),
    .Q(\digitop_pav2.sec_inst.reg160[52] ));
 dfrtp_1 _23672_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00629_),
    .RESET_B(net997),
    .Q(\digitop_pav2.sec_inst.reg160[53] ));
 dfrtp_1 _23673_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00630_),
    .RESET_B(net997),
    .Q(\digitop_pav2.sec_inst.reg160[54] ));
 dfrtp_1 _23674_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00631_),
    .RESET_B(net999),
    .Q(\digitop_pav2.sec_inst.reg160[55] ));
 dfrtp_1 _23675_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00632_),
    .RESET_B(net999),
    .Q(\digitop_pav2.sec_inst.reg160[56] ));
 dfrtp_1 _23676_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00633_),
    .RESET_B(net999),
    .Q(\digitop_pav2.sec_inst.reg160[57] ));
 dfrtp_1 _23677_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00634_),
    .RESET_B(net999),
    .Q(\digitop_pav2.sec_inst.reg160[58] ));
 dfrtp_1 _23678_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00635_),
    .RESET_B(net998),
    .Q(\digitop_pav2.sec_inst.reg160[59] ));
 dfrtp_1 _23679_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00636_),
    .RESET_B(net999),
    .Q(\digitop_pav2.sec_inst.reg160[60] ));
 dfrtp_1 _23680_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00637_),
    .RESET_B(net998),
    .Q(\digitop_pav2.sec_inst.reg160[61] ));
 dfrtp_1 _23681_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00638_),
    .RESET_B(net998),
    .Q(\digitop_pav2.sec_inst.reg160[62] ));
 dfrtp_1 _23682_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00639_),
    .RESET_B(net997),
    .Q(\digitop_pav2.sec_inst.reg160[63] ));
 dfstp_1 _23683_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00640_),
    .SET_B(net1003),
    .Q(\digitop_pav2.sec_inst.shift_in.s12.q[0] ));
 dfrtp_1 _23684_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00641_),
    .RESET_B(net1002),
    .Q(\digitop_pav2.sec_inst.shift_in.s12.q[1] ));
 dfrtp_1 _23685_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00642_),
    .RESET_B(net1002),
    .Q(\digitop_pav2.sec_inst.shift_in.s12.q[2] ));
 dfrtp_1 _23686_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00643_),
    .RESET_B(net1002),
    .Q(\digitop_pav2.sec_inst.shift_in.s12.q[3] ));
 dfrtp_1 _23687_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00644_),
    .RESET_B(net1003),
    .Q(\digitop_pav2.sec_inst.shift_in.s12.q[4] ));
 dfrtp_1 _23688_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00645_),
    .RESET_B(net1003),
    .Q(\digitop_pav2.sec_inst.shift_in.s12.q[5] ));
 dfrtp_1 _23689_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00646_),
    .RESET_B(net1003),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[6] ));
 dfrtp_1 _23690_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00647_),
    .RESET_B(net1003),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[7] ));
 dfstp_1 _23691_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00648_),
    .SET_B(net982),
    .Q(\digitop_pav2.sec_inst.shift_in.s11.q[0] ));
 dfrtp_1 _23692_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00649_),
    .RESET_B(net985),
    .Q(\digitop_pav2.sec_inst.shift_in.s11.q[1] ));
 dfrtp_1 _23693_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00650_),
    .RESET_B(net985),
    .Q(\digitop_pav2.sec_inst.shift_in.s11.q[2] ));
 dfrtp_1 _23694_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00651_),
    .RESET_B(net982),
    .Q(\digitop_pav2.sec_inst.shift_in.s11.q[3] ));
 dfrtp_1 _23695_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00652_),
    .RESET_B(net982),
    .Q(\digitop_pav2.sec_inst.shift_in.s11.q[4] ));
 dfrtp_1 _23696_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00653_),
    .RESET_B(net983),
    .Q(\digitop_pav2.sec_inst.shift_in.s11.q[5] ));
 dfrtp_1 _23697_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00654_),
    .RESET_B(net982),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[14] ));
 dfrtp_1 _23698_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00655_),
    .RESET_B(net991),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[15] ));
 dfstp_1 _23699_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00656_),
    .SET_B(net1004),
    .Q(\digitop_pav2.sec_inst.shift_in.s10.q[0] ));
 dfrtp_1 _23700_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00657_),
    .RESET_B(net1004),
    .Q(\digitop_pav2.sec_inst.shift_in.s10.q[1] ));
 dfrtp_1 _23701_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00658_),
    .RESET_B(net1004),
    .Q(\digitop_pav2.sec_inst.shift_in.s10.q[2] ));
 dfrtp_1 _23702_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00659_),
    .RESET_B(net1004),
    .Q(\digitop_pav2.sec_inst.shift_in.s10.q[3] ));
 dfrtp_1 _23703_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00660_),
    .RESET_B(net1002),
    .Q(\digitop_pav2.sec_inst.shift_in.s10.q[4] ));
 dfrtp_1 _23704_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00661_),
    .RESET_B(net1002),
    .Q(\digitop_pav2.sec_inst.shift_in.s10.q[5] ));
 dfrtp_1 _23705_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00662_),
    .RESET_B(net1004),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[22] ));
 dfrtp_1 _23706_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00663_),
    .RESET_B(net1002),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[23] ));
 dfstp_1 _23707_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00664_),
    .SET_B(net989),
    .Q(\digitop_pav2.sec_inst.shift_in.s1.q[0] ));
 dfrtp_1 _23708_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00665_),
    .RESET_B(net987),
    .Q(\digitop_pav2.sec_inst.shift_in.s1.q[1] ));
 dfrtp_1 _23709_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00666_),
    .RESET_B(net980),
    .Q(\digitop_pav2.sec_inst.shift_in.s1.q[2] ));
 dfrtp_1 _23710_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00667_),
    .RESET_B(net980),
    .Q(\digitop_pav2.sec_inst.shift_in.s1.q[3] ));
 dfrtp_1 _23711_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00668_),
    .RESET_B(net980),
    .Q(\digitop_pav2.sec_inst.shift_in.s1.q[4] ));
 dfrtp_1 _23712_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00669_),
    .RESET_B(net980),
    .Q(\digitop_pav2.sec_inst.shift_in.s1.q[5] ));
 dfrtp_1 _23713_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00670_),
    .RESET_B(net980),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[94] ));
 dfrtp_1 _23714_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00671_),
    .RESET_B(net992),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[95] ));
 dfstp_1 _23715_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00672_),
    .SET_B(net985),
    .Q(\digitop_pav2.sec_inst.shift_in.s8.q[0] ));
 dfrtp_1 _23716_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00673_),
    .RESET_B(net985),
    .Q(\digitop_pav2.sec_inst.shift_in.s8.q[1] ));
 dfrtp_1 _23717_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00674_),
    .RESET_B(net985),
    .Q(\digitop_pav2.sec_inst.shift_in.s8.q[2] ));
 dfrtp_1 _23718_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00675_),
    .RESET_B(net985),
    .Q(\digitop_pav2.sec_inst.shift_in.s8.q[3] ));
 dfrtp_1 _23719_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00676_),
    .RESET_B(net1003),
    .Q(\digitop_pav2.sec_inst.shift_in.s8.q[4] ));
 dfrtp_1 _23720_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00677_),
    .RESET_B(net1003),
    .Q(\digitop_pav2.sec_inst.shift_in.s8.q[5] ));
 dfrtp_1 _23721_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00678_),
    .RESET_B(net991),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[38] ));
 dfrtp_1 _23722_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00679_),
    .RESET_B(net991),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[39] ));
 dfstp_1 _23723_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(net1642),
    .SET_B(net982),
    .Q(\digitop_pav2.sec_inst.shift_in.s7.q[0] ));
 dfrtp_1 _23724_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00681_),
    .RESET_B(net981),
    .Q(\digitop_pav2.sec_inst.shift_in.s7.q[1] ));
 dfrtp_1 _23725_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00682_),
    .RESET_B(net980),
    .Q(\digitop_pav2.sec_inst.shift_in.s7.q[2] ));
 dfrtp_1 _23726_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00683_),
    .RESET_B(net981),
    .Q(\digitop_pav2.sec_inst.shift_in.s7.q[3] ));
 dfrtp_1 _23727_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00684_),
    .RESET_B(net981),
    .Q(\digitop_pav2.sec_inst.shift_in.s7.q[4] ));
 dfrtp_1 _23728_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00685_),
    .RESET_B(net981),
    .Q(\digitop_pav2.sec_inst.shift_in.s7.q[5] ));
 dfrtp_1 _23729_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00686_),
    .RESET_B(net981),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[46] ));
 dfrtp_1 _23730_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00687_),
    .RESET_B(net983),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[47] ));
 dfstp_1 _23731_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00688_),
    .SET_B(net992),
    .Q(\digitop_pav2.sec_inst.shift_in.s6.q[0] ));
 dfrtp_1 _23732_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00689_),
    .RESET_B(net991),
    .Q(\digitop_pav2.sec_inst.shift_in.s6.q[1] ));
 dfrtp_1 _23733_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00690_),
    .RESET_B(net1004),
    .Q(\digitop_pav2.sec_inst.shift_in.s6.q[2] ));
 dfrtp_1 _23734_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00691_),
    .RESET_B(net1002),
    .Q(\digitop_pav2.sec_inst.shift_in.s6.q[3] ));
 dfrtp_1 _23735_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00692_),
    .RESET_B(net1002),
    .Q(\digitop_pav2.sec_inst.shift_in.s6.q[4] ));
 dfrtp_1 _23736_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00693_),
    .RESET_B(net1002),
    .Q(\digitop_pav2.sec_inst.shift_in.s6.q[5] ));
 dfrtp_1 _23737_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00694_),
    .RESET_B(net1003),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[54] ));
 dfrtp_1 _23738_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00695_),
    .RESET_B(net991),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[55] ));
 dfstp_1 _23739_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00696_),
    .SET_B(net987),
    .Q(\digitop_pav2.sec_inst.shift_in.s5.q[0] ));
 dfrtp_1 _23740_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00697_),
    .RESET_B(net990),
    .Q(\digitop_pav2.sec_inst.shift_in.s5.q[1] ));
 dfrtp_1 _23741_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00698_),
    .RESET_B(net987),
    .Q(\digitop_pav2.sec_inst.shift_in.s5.q[2] ));
 dfrtp_1 _23742_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00699_),
    .RESET_B(net980),
    .Q(\digitop_pav2.sec_inst.shift_in.s5.q[3] ));
 dfrtp_1 _23743_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00700_),
    .RESET_B(net980),
    .Q(\digitop_pav2.sec_inst.shift_in.s5.q[4] ));
 dfrtp_1 _23744_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00701_),
    .RESET_B(net980),
    .Q(\digitop_pav2.sec_inst.shift_in.s5.q[5] ));
 dfrtp_1 _23745_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00702_),
    .RESET_B(net980),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[62] ));
 dfrtp_1 _23746_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00703_),
    .RESET_B(net991),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[63] ));
 dfstp_1 _23747_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00704_),
    .SET_B(net997),
    .Q(\digitop_pav2.sec_inst.shift_in.s4.q[0] ));
 dfrtp_1 _23748_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00705_),
    .RESET_B(net1000),
    .Q(\digitop_pav2.sec_inst.shift_in.s4.q[1] ));
 dfrtp_1 _23749_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00706_),
    .RESET_B(net1000),
    .Q(\digitop_pav2.sec_inst.shift_in.s4.q[2] ));
 dfrtp_1 _23750_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00707_),
    .RESET_B(net1000),
    .Q(\digitop_pav2.sec_inst.shift_in.s4.q[3] ));
 dfrtp_1 _23751_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00708_),
    .RESET_B(net1004),
    .Q(\digitop_pav2.sec_inst.shift_in.s4.q[4] ));
 dfrtp_1 _23752_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00709_),
    .RESET_B(net997),
    .Q(\digitop_pav2.sec_inst.shift_in.s4.q[5] ));
 dfrtp_1 _23753_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00710_),
    .RESET_B(net1004),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[70] ));
 dfrtp_1 _23754_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00711_),
    .RESET_B(net992),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[71] ));
 dfstp_1 _23755_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00712_),
    .SET_B(net991),
    .Q(\digitop_pav2.sec_inst.shift_in.s3.q[0] ));
 dfrtp_1 _23756_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00713_),
    .RESET_B(net987),
    .Q(\digitop_pav2.sec_inst.shift_in.s3.q[1] ));
 dfrtp_1 _23757_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00714_),
    .RESET_B(net987),
    .Q(\digitop_pav2.sec_inst.shift_in.s3.q[2] ));
 dfrtp_1 _23758_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00715_),
    .RESET_B(net987),
    .Q(\digitop_pav2.sec_inst.shift_in.s3.q[3] ));
 dfrtp_1 _23759_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00716_),
    .RESET_B(net987),
    .Q(\digitop_pav2.sec_inst.shift_in.s3.q[4] ));
 dfrtp_1 _23760_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00717_),
    .RESET_B(net988),
    .Q(\digitop_pav2.sec_inst.shift_in.s3.q[5] ));
 dfrtp_1 _23761_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00718_),
    .RESET_B(net989),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[78] ));
 dfrtp_1 _23762_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00719_),
    .RESET_B(net991),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[79] ));
 dfstp_1 _23763_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00720_),
    .SET_B(net992),
    .Q(\digitop_pav2.sec_inst.shift_in.s2.q[0] ));
 dfrtp_1 _23764_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00721_),
    .RESET_B(net997),
    .Q(\digitop_pav2.sec_inst.shift_in.s2.q[1] ));
 dfrtp_1 _23765_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00722_),
    .RESET_B(net1000),
    .Q(\digitop_pav2.sec_inst.shift_in.s2.q[2] ));
 dfrtp_1 _23766_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00723_),
    .RESET_B(net991),
    .Q(\digitop_pav2.sec_inst.shift_in.s2.q[3] ));
 dfrtp_1 _23767_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00724_),
    .RESET_B(net992),
    .Q(\digitop_pav2.sec_inst.shift_in.s2.q[4] ));
 dfrtp_1 _23768_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00725_),
    .RESET_B(net992),
    .Q(\digitop_pav2.sec_inst.shift_in.s2.q[5] ));
 dfrtp_1 _23769_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00726_),
    .RESET_B(net1002),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[86] ));
 dfrtp_1 _23770_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00727_),
    .RESET_B(net992),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[87] ));
 dfstp_1 _23771_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00728_),
    .SET_B(net989),
    .Q(\digitop_pav2.sec_inst.reg160[0] ));
 dfrtp_1 _23772_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00729_),
    .RESET_B(net988),
    .Q(\digitop_pav2.sec_inst.reg160[1] ));
 dfrtp_1 _23773_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00730_),
    .RESET_B(net988),
    .Q(\digitop_pav2.sec_inst.reg160[2] ));
 dfrtp_1 _23774_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00731_),
    .RESET_B(net987),
    .Q(\digitop_pav2.sec_inst.reg160[3] ));
 dfrtp_1 _23775_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00732_),
    .RESET_B(net987),
    .Q(\digitop_pav2.sec_inst.reg160[4] ));
 dfrtp_1 _23776_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00733_),
    .RESET_B(net988),
    .Q(\digitop_pav2.sec_inst.reg160[5] ));
 dfrtp_1 _23777_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00734_),
    .RESET_B(net988),
    .Q(\digitop_pav2.sec_inst.reg160[6] ));
 dfrtp_1 _23778_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00735_),
    .RESET_B(net988),
    .Q(\digitop_pav2.sec_inst.reg160[7] ));
 dfrtp_1 _23779_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00736_),
    .RESET_B(net988),
    .Q(\digitop_pav2.sec_inst.reg160[8] ));
 dfrtp_1 _23780_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00737_),
    .RESET_B(net988),
    .Q(\digitop_pav2.sec_inst.reg160[9] ));
 dfrtp_1 _23781_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00738_),
    .RESET_B(net988),
    .Q(\digitop_pav2.sec_inst.reg160[10] ));
 dfrtp_1 _23782_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00739_),
    .RESET_B(net988),
    .Q(\digitop_pav2.sec_inst.reg160[11] ));
 dfrtp_1 _23783_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00740_),
    .RESET_B(net989),
    .Q(\digitop_pav2.sec_inst.reg160[12] ));
 dfrtp_1 _23784_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00741_),
    .RESET_B(net989),
    .Q(\digitop_pav2.sec_inst.reg160[13] ));
 dfrtp_1 _23785_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00742_),
    .RESET_B(net993),
    .Q(\digitop_pav2.sec_inst.reg160[14] ));
 dfrtp_1 _23786_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00743_),
    .RESET_B(net992),
    .Q(\digitop_pav2.sec_inst.reg160[15] ));
 dfrtp_2 _23787_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00744_),
    .RESET_B(net989),
    .Q(\digitop_pav2.sec_inst.shift_in.st[0] ));
 dfrtp_1 _23788_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00745_),
    .RESET_B(net989),
    .Q(\digitop_pav2.sec_inst.shift_in.st[1] ));
 dfrtp_2 _23789_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00746_),
    .RESET_B(net990),
    .Q(\digitop_pav2.sec_inst.shift_in.st[2] ));
 dfrtp_1 _23790_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00747_),
    .RESET_B(net987),
    .Q(\digitop_pav2.sec_inst.shift_in.st[3] ));
 dfrtp_1 _23791_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00748_),
    .RESET_B(net989),
    .Q(\digitop_pav2.sec_inst.shift_in.st[4] ));
 dfxtp_1 _23792_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00749_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[0] ));
 dfxtp_1 _23793_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00750_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[1] ));
 dfxtp_1 _23794_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00751_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[2] ));
 dfxtp_1 _23795_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00752_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[3] ));
 dfxtp_1 _23796_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00753_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[4] ));
 dfxtp_1 _23797_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00754_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[5] ));
 dfxtp_1 _23798_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00755_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[6] ));
 dfxtp_1 _23799_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00756_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[7] ));
 dfxtp_1 _23800_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00757_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[8] ));
 dfxtp_1 _23801_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00758_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[9] ));
 dfxtp_1 _23802_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00759_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[10] ));
 dfxtp_1 _23803_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00760_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[11] ));
 dfxtp_1 _23804_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00761_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[12] ));
 dfxtp_1 _23805_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00762_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[13] ));
 dfxtp_1 _23806_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00763_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[14] ));
 dfxtp_1 _23807_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00764_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[15] ));
 dfxtp_1 _23808_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00765_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[16] ));
 dfxtp_1 _23809_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00766_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[17] ));
 dfxtp_1 _23810_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00767_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[18] ));
 dfxtp_1 _23811_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00768_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[19] ));
 dfxtp_1 _23812_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00769_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[20] ));
 dfxtp_1 _23813_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00770_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[21] ));
 dfxtp_1 _23814_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00771_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[22] ));
 dfxtp_1 _23815_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00772_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[23] ));
 dfxtp_1 _23816_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00773_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[24] ));
 dfxtp_1 _23817_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00774_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[25] ));
 dfxtp_1 _23818_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00775_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[26] ));
 dfxtp_1 _23819_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00776_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[27] ));
 dfxtp_1 _23820_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00777_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[28] ));
 dfxtp_1 _23821_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00778_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[29] ));
 dfxtp_1 _23822_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00779_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[30] ));
 dfxtp_1 _23823_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00780_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[31] ));
 dfxtp_1 _23824_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00781_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[32] ));
 dfxtp_1 _23825_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00782_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[33] ));
 dfxtp_1 _23826_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00783_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[34] ));
 dfxtp_1 _23827_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00784_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[35] ));
 dfxtp_1 _23828_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00785_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[36] ));
 dfxtp_1 _23829_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00786_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[37] ));
 dfxtp_1 _23830_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00787_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[38] ));
 dfxtp_1 _23831_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00788_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[39] ));
 dfxtp_1 _23832_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00789_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[40] ));
 dfxtp_1 _23833_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00790_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[41] ));
 dfxtp_1 _23834_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00791_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[42] ));
 dfxtp_1 _23835_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00792_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[43] ));
 dfxtp_1 _23836_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00793_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[44] ));
 dfxtp_1 _23837_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00794_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[45] ));
 dfxtp_1 _23838_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00795_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[46] ));
 dfxtp_1 _23839_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00796_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[47] ));
 dfxtp_1 _23840_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00797_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[48] ));
 dfxtp_1 _23841_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00798_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[49] ));
 dfxtp_1 _23842_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00799_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[50] ));
 dfxtp_1 _23843_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00800_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[51] ));
 dfxtp_1 _23844_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00801_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[52] ));
 dfxtp_1 _23845_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00802_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[53] ));
 dfxtp_1 _23846_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00803_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[54] ));
 dfxtp_1 _23847_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00804_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[55] ));
 dfxtp_1 _23848_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00805_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[56] ));
 dfxtp_1 _23849_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00806_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[57] ));
 dfxtp_1 _23850_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00807_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[58] ));
 dfxtp_1 _23851_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00808_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[59] ));
 dfxtp_1 _23852_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00809_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[60] ));
 dfxtp_1 _23853_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00810_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[61] ));
 dfxtp_1 _23854_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00811_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[62] ));
 dfxtp_1 _23855_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00812_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[63] ));
 dfxtp_1 _23856_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00813_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[64] ));
 dfxtp_1 _23857_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00814_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[65] ));
 dfxtp_1 _23858_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00815_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[66] ));
 dfxtp_1 _23859_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00816_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[67] ));
 dfxtp_1 _23860_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00817_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[68] ));
 dfxtp_1 _23861_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00818_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[69] ));
 dfxtp_1 _23862_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00819_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[70] ));
 dfxtp_1 _23863_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00820_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[71] ));
 dfxtp_1 _23864_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00821_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[72] ));
 dfxtp_1 _23865_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00822_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[73] ));
 dfxtp_1 _23866_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00823_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[74] ));
 dfxtp_1 _23867_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00824_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[75] ));
 dfxtp_1 _23868_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00825_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[76] ));
 dfxtp_1 _23869_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00826_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[77] ));
 dfxtp_1 _23870_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00827_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[78] ));
 dfxtp_1 _23871_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00828_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[79] ));
 dfxtp_1 _23872_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00829_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[80] ));
 dfxtp_1 _23873_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00830_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[81] ));
 dfxtp_1 _23874_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00831_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[82] ));
 dfxtp_1 _23875_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00832_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[83] ));
 dfxtp_1 _23876_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00833_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[84] ));
 dfxtp_1 _23877_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00834_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[85] ));
 dfxtp_1 _23878_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00835_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[86] ));
 dfxtp_1 _23879_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00836_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[87] ));
 dfxtp_1 _23880_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00837_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[88] ));
 dfxtp_1 _23881_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00838_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[89] ));
 dfxtp_1 _23882_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00839_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[90] ));
 dfxtp_1 _23883_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00840_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[91] ));
 dfxtp_1 _23884_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00841_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[92] ));
 dfxtp_1 _23885_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00842_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[93] ));
 dfxtp_1 _23886_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00843_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[94] ));
 dfxtp_1 _23887_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00844_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[95] ));
 dfxtp_1 _23888_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00845_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[96] ));
 dfxtp_1 _23889_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00846_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[97] ));
 dfxtp_1 _23890_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00847_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[98] ));
 dfxtp_1 _23891_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00848_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[99] ));
 dfxtp_1 _23892_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00849_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[100] ));
 dfxtp_1 _23893_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00850_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[101] ));
 dfxtp_1 _23894_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00851_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[102] ));
 dfxtp_1 _23895_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00852_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[103] ));
 dfxtp_1 _23896_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00853_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[104] ));
 dfxtp_1 _23897_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00854_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[105] ));
 dfxtp_1 _23898_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00855_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[106] ));
 dfxtp_1 _23899_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00856_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[107] ));
 dfxtp_1 _23900_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00857_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[108] ));
 dfxtp_1 _23901_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00858_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[109] ));
 dfxtp_1 _23902_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00859_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[110] ));
 dfxtp_1 _23903_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00860_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[111] ));
 dfxtp_1 _23904_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00861_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[112] ));
 dfxtp_1 _23905_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00862_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[113] ));
 dfxtp_1 _23906_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00863_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[114] ));
 dfxtp_1 _23907_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00864_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[115] ));
 dfxtp_1 _23908_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00865_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[116] ));
 dfxtp_1 _23909_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00866_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[117] ));
 dfxtp_1 _23910_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00867_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[118] ));
 dfxtp_1 _23911_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00868_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[119] ));
 dfxtp_1 _23912_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00869_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[120] ));
 dfxtp_1 _23913_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00870_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[121] ));
 dfxtp_1 _23914_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00871_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[122] ));
 dfxtp_1 _23915_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00872_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[123] ));
 dfxtp_1 _23916_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00873_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[124] ));
 dfxtp_1 _23917_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00874_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[125] ));
 dfxtp_1 _23918_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00875_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[126] ));
 dfxtp_1 _23919_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00876_),
    .Q(\digitop_pav2.sec_inst.r128.reg128_o[127] ));
 dfrtp_1 _23920_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00877_),
    .RESET_B(net984),
    .Q(\digitop_pav2.sec_inst.shift_out.j_ctr[0] ));
 dfrtp_1 _23921_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00878_),
    .RESET_B(net984),
    .Q(\digitop_pav2.sec_inst.shift_out.j_ctr[1] ));
 dfrtp_1 _23922_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00879_),
    .RESET_B(net984),
    .Q(\digitop_pav2.sec_inst.shift_out.j_ctr[2] ));
 dfrtp_1 _23923_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00880_),
    .RESET_B(net984),
    .Q(\digitop_pav2.sec_inst.shift_out.j_ctr[3] ));
 dfrtp_1 _23924_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00881_),
    .RESET_B(net984),
    .Q(\digitop_pav2.sec_inst.shift_out.j_ctr[4] ));
 dfrtp_1 _23925_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00882_),
    .RESET_B(net984),
    .Q(\digitop_pav2.sec_inst.shift_out.j_ctr[5] ));
 dfrtp_4 _23926_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00883_),
    .RESET_B(net984),
    .Q(\digitop_pav2.sec_inst.shift_out.j_ctr[6] ));
 dfstp_1 _23927_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00884_),
    .SET_B(net983),
    .Q(\digitop_pav2.sec_inst.shift_in.s9.q[0] ));
 dfrtp_1 _23928_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00885_),
    .RESET_B(net983),
    .Q(\digitop_pav2.sec_inst.shift_in.s9.q[1] ));
 dfrtp_1 _23929_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00886_),
    .RESET_B(net982),
    .Q(\digitop_pav2.sec_inst.shift_in.s9.q[2] ));
 dfrtp_1 _23930_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00887_),
    .RESET_B(net982),
    .Q(\digitop_pav2.sec_inst.shift_in.s9.q[3] ));
 dfrtp_1 _23931_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00888_),
    .RESET_B(net982),
    .Q(\digitop_pav2.sec_inst.shift_in.s9.q[4] ));
 dfrtp_1 _23932_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00889_),
    .RESET_B(net982),
    .Q(\digitop_pav2.sec_inst.shift_in.s9.q[5] ));
 dfrtp_1 _23933_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00890_),
    .RESET_B(net982),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[30] ));
 dfrtp_1 _23934_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00891_),
    .RESET_B(net991),
    .Q(\digitop_pav2.sec_inst.ld_r.reg96_i[31] ));
 dfrtp_2 _23935_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00892_),
    .RESET_B(net986),
    .Q(\digitop_pav2.sec_inst.shift_out.ctr[0] ));
 dfrtp_2 _23936_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00893_),
    .RESET_B(net986),
    .Q(\digitop_pav2.sec_inst.shift_out.ctr[1] ));
 dfrtp_1 _23937_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00894_),
    .RESET_B(net984),
    .Q(\digitop_pav2.sec_inst.shift_out.ctr[2] ));
 dfrtp_1 _23938_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_00895_),
    .RESET_B(net984),
    .Q(\digitop_pav2.sec_inst.shift_out.ctr[3] ));
 dfrtp_1 _23939_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(net1654),
    .RESET_B(net1006),
    .Q(\digitop_pav2.sec_inst.ld_mem.round_i ));
 dfstp_1 _23940_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00064_),
    .SET_B(net1269),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.state[0] ));
 dfrtp_1 _23941_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00069_),
    .RESET_B(net1268),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.state[1] ));
 dfrtp_1 _23942_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00070_),
    .RESET_B(net1268),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.state[2] ));
 dfrtp_1 _23943_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00071_),
    .RESET_B(net1269),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.select_valid_o ));
 dfrtp_2 _23944_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00072_),
    .RESET_B(net1269),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.state[4] ));
 dfrtp_1 _23945_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00073_),
    .RESET_B(net1268),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.state[5] ));
 dfrtp_2 _23946_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00074_),
    .RESET_B(net1268),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.state[6] ));
 dfrtp_1 _23947_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00075_),
    .RESET_B(net1268),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.state[7] ));
 dfrtp_2 _23948_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00076_),
    .RESET_B(net1269),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.r_invent2_o ));
 dfrtp_1 _23949_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00077_),
    .RESET_B(net1268),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.state[9] ));
 dfrtp_1 _23950_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00065_),
    .RESET_B(net1269),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.state[10] ));
 dfrtp_1 _23951_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00066_),
    .RESET_B(net1268),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.state[11] ));
 dfrtp_2 _23952_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00067_),
    .RESET_B(net1268),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.state[12] ));
 dfrtp_1 _23953_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00068_),
    .RESET_B(net1269),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.r_invent3_o ));
 dfxtp_1 _23954_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00897_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[6] ));
 dfxtp_1 _23955_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00898_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.rcon_i[7] ));
 dfxtp_1 _23956_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00899_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[0] ));
 dfxtp_1 _23957_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00900_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[1] ));
 dfxtp_1 _23958_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00901_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[2] ));
 dfxtp_1 _23959_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00902_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[3] ));
 dfxtp_1 _23960_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00903_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[4] ));
 dfxtp_1 _23961_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00904_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[5] ));
 dfxtp_1 _23962_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00905_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[6] ));
 dfxtp_1 _23963_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00906_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[7] ));
 dfxtp_1 _23964_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00907_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[8] ));
 dfxtp_1 _23965_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00908_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[9] ));
 dfxtp_1 _23966_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00909_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[10] ));
 dfxtp_1 _23967_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00910_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[11] ));
 dfxtp_1 _23968_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00911_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[12] ));
 dfxtp_1 _23969_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00912_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[13] ));
 dfxtp_1 _23970_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00913_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[14] ));
 dfxtp_1 _23971_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00914_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf2[15] ));
 dfrtp_1 _23972_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00915_),
    .RESET_B(net1816),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[0] ));
 dfrtp_1 _23973_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00916_),
    .RESET_B(net1250),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[1] ));
 dfrtp_1 _23974_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00917_),
    .RESET_B(net1816),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[2] ));
 dfrtp_1 _23975_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00918_),
    .RESET_B(net1816),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[3] ));
 dfrtp_1 _23976_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00919_),
    .RESET_B(net1250),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr1[4] ));
 dfxtp_1 _23977_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00920_),
    .Q(\digitop_pav2.func_rng_data[0] ));
 dfxtp_1 _23978_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00921_),
    .Q(\digitop_pav2.func_rng_data[1] ));
 dfxtp_1 _23979_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00922_),
    .Q(\digitop_pav2.func_rng_data[2] ));
 dfxtp_1 _23980_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00923_),
    .Q(\digitop_pav2.func_rng_data[3] ));
 dfxtp_1 _23981_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00924_),
    .Q(\digitop_pav2.func_rng_data[4] ));
 dfxtp_1 _23982_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00925_),
    .Q(\digitop_pav2.func_rng_data[5] ));
 dfxtp_1 _23983_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00926_),
    .Q(\digitop_pav2.func_rng_data[6] ));
 dfxtp_2 _23984_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00927_),
    .Q(\digitop_pav2.func_rng_data[7] ));
 dfxtp_2 _23985_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00928_),
    .Q(\digitop_pav2.func_rng_data[8] ));
 dfxtp_2 _23986_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00929_),
    .Q(\digitop_pav2.func_rng_data[9] ));
 dfxtp_1 _23987_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00930_),
    .Q(\digitop_pav2.func_rng_data[10] ));
 dfxtp_1 _23988_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00931_),
    .Q(\digitop_pav2.func_rng_data[11] ));
 dfxtp_1 _23989_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00932_),
    .Q(\digitop_pav2.func_rng_data[12] ));
 dfxtp_1 _23990_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00933_),
    .Q(\digitop_pav2.func_rng_data[13] ));
 dfxtp_1 _23991_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00934_),
    .Q(\digitop_pav2.func_rng_data[14] ));
 dfxtp_1 _23992_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(_00935_),
    .Q(\digitop_pav2.func_rng_data[15] ));
 dfxtp_1 _23993_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(\digitop_pav2.rng_inst.rng_trngx_pav2.ff1 ),
    .Q(\digitop_pav2.rng_inst.rng_prngx_pav2.trngx_data_i ));
 dfxtp_1 _23994_ (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(\digitop_pav2.rng_inst.rng_trngx_pav2.xor_data ),
    .Q(\digitop_pav2.rng_inst.rng_trngx_pav2.ff1 ));
 dfrtp_2 _23995_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00936_),
    .RESET_B(net1450),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.en_i ));
 dfrtp_1 _23996_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00937_),
    .RESET_B(net1223),
    .Q(\digitop_pav2.g_reqrn ));
 dfrtp_1 _23997_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00938_),
    .RESET_B(net1223),
    .Q(\digitop_pav2.g_queryrep ));
 dfrtp_1 _23998_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00939_),
    .RESET_B(net1223),
    .Q(\digitop_pav2.g_queryadj ));
 dfrtp_1 _23999_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00940_),
    .RESET_B(net1223),
    .Q(\digitop_pav2.access_inst.access_check0.g_write_i ));
 dfrtp_1 _24000_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00941_),
    .RESET_B(net1223),
    .Q(\digitop_pav2.g_query ));
 dfrtp_1 _24001_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00942_),
    .RESET_B(net1223),
    .Q(\digitop_pav2.g_select ));
 dfrtp_1 _24002_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00943_),
    .RESET_B(net1224),
    .Q(\digitop_pav2.ack_inst.g_ack_i ));
 dfrtp_1 _24003_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_00944_),
    .RESET_B(net1455),
    .Q(\digitop_pav2.pie_inst.fsm.comp_tari_ff ));
 dfrtp_4 _24004_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00945_),
    .RESET_B(net1223),
    .Q(\digitop_pav2.access_inst.access_check0.g_propwrite_i ));
 dfrtp_1 _24005_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00946_),
    .RESET_B(net1224),
    .Q(\digitop_pav2.access_inst.access_check0.g_read_i ));
 dfrtp_1 _24006_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00947_),
    .RESET_B(net1223),
    .Q(\digitop_pav2.access_inst.access_check0.g_activate_i ));
 dfrtp_1 _24007_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00948_),
    .RESET_B(net1223),
    .Q(\digitop_pav2.proc_ctrl_inst.cmd.g_sec_auth_o ));
 dfrtp_1 _24008_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00949_),
    .RESET_B(net973),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.invalid ));
 dfrtp_1 _24009_ (.CLK(\digitop_pav2.clkx_irreg_clk ),
    .D(net1611),
    .RESET_B(_00214_),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.t2.jalido ));
 dfrtp_4 _24010_ (.CLK(_00216_),
    .D(_00145_),
    .RESET_B(_00215_),
    .Q(\digitop_pav2.proc_ctrl_inst.int_timeout_t2 ));
 dfrtp_1 _24011_ (.CLK(\digitop_pav2.fm0x_clk_for_proc_ctrl ),
    .D(_00950_),
    .RESET_B(_00217_),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[0] ));
 dfrtp_1 _24012_ (.CLK(\digitop_pav2.fm0x_clk_for_proc_ctrl ),
    .D(_00951_),
    .RESET_B(_00218_),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[1] ));
 dfrtp_1 _24013_ (.CLK(\digitop_pav2.fm0x_clk_for_proc_ctrl ),
    .D(_00952_),
    .RESET_B(_00219_),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[2] ));
 dfrtp_1 _24014_ (.CLK(\digitop_pav2.fm0x_clk_for_proc_ctrl ),
    .D(_00953_),
    .RESET_B(_00220_),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[3] ));
 dfrtp_1 _24015_ (.CLK(\digitop_pav2.fm0x_clk_for_proc_ctrl ),
    .D(_00954_),
    .RESET_B(_00221_),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.ctr.ctr2[4] ));
 dfrtp_1 _24016_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00955_),
    .RESET_B(net1449),
    .Q(\digitop_pav2.proc_ctrl_inst.profsm.r1_rise_ff ));
 dfrtp_4 _24017_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(\digitop_pav2.proc_ctrl_inst.cmdfsm.n_pass_t1_i ),
    .RESET_B(net1250),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.pass_t1_i ));
 dfrtp_1 _24018_ (.CLK(\digitop_pav2.fm0x_clk_for_proc_ctrl ),
    .D(_00144_),
    .RESET_B(_00222_),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.ctr.pass_t2 ));
 dfrtp_1 _24019_ (.CLK(\digitop_pav2.fm0x_clk_for_proc_ctrl ),
    .D(_00956_),
    .RESET_B(_00223_),
    .Q(\digitop_pav2.proc_ctrl_inst.timeout.ctr.pass_t2_flag ));
 dfrtp_1 _24020_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00957_),
    .RESET_B(net1224),
    .Q(\digitop_pav2.proc_ctrl_inst.cmd.state[0] ));
 dfrtp_1 _24021_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00958_),
    .RESET_B(net1224),
    .Q(\digitop_pav2.proc_ctrl_inst.cmd.state[1] ));
 dfrtp_4 _24022_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00959_),
    .RESET_B(net1224),
    .Q(\digitop_pav2.proc_ctrl_inst.cmd.state[2] ));
 dfrtp_4 _24023_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00960_),
    .RESET_B(net1224),
    .Q(\digitop_pav2.proc_ctrl_inst.cmd.state[3] ));
 dfrtp_1 _24024_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00961_),
    .RESET_B(net1223),
    .Q(\digitop_pav2.proc_ctrl_inst.cmd.state[4] ));
 dfrtp_4 _24025_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00962_),
    .RESET_B(net1224),
    .Q(\digitop_pav2.proc_ctrl_inst.cmd.state[5] ));
 dfstp_1 _24026_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00963_),
    .SET_B(_00224_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[0] ));
 dfstp_1 _24027_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00964_),
    .SET_B(_00225_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[1] ));
 dfstp_1 _24028_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00965_),
    .SET_B(_00226_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[2] ));
 dfstp_1 _24029_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00966_),
    .SET_B(_00227_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[3] ));
 dfstp_1 _24030_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00967_),
    .SET_B(_00228_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[4] ));
 dfstp_1 _24031_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00968_),
    .SET_B(_00229_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[5] ));
 dfstp_1 _24032_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00969_),
    .SET_B(_00230_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[6] ));
 dfstp_1 _24033_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00970_),
    .SET_B(_00231_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.ctr[7] ));
 dfrtp_1 _24034_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00971_),
    .RESET_B(_00232_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.cmdctr_end3 ));
 dfrtp_1 _24035_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00972_),
    .RESET_B(_00233_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.par1_en_ff ));
 dfrtp_1 _24036_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00973_),
    .RESET_B(_00234_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.par2_en_ff ));
 dfrtp_1 _24037_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00974_),
    .RESET_B(_00235_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.par3_en_ff ));
 dfxtp_1 _24038_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00975_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[0] ));
 dfxtp_1 _24039_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00976_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[1] ));
 dfxtp_1 _24040_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00977_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[2] ));
 dfxtp_1 _24041_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00978_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[3] ));
 dfxtp_1 _24042_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00979_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[4] ));
 dfxtp_1 _24043_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00980_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[5] ));
 dfxtp_1 _24044_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00981_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[6] ));
 dfxtp_1 _24045_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00982_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[7] ));
 dfxtp_1 _24046_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00983_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[8] ));
 dfxtp_1 _24047_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00984_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[9] ));
 dfxtp_1 _24048_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00985_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[10] ));
 dfxtp_1 _24049_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00986_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[11] ));
 dfxtp_1 _24050_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00987_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[12] ));
 dfxtp_1 _24051_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00988_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[13] ));
 dfxtp_1 _24052_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00989_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[14] ));
 dfxtp_1 _24053_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00990_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.handle_i[15] ));
 dfrtp_2 _24054_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(net475),
    .RESET_B(net1225),
    .Q(\digitop_pav2.pie_inst.fsm.state[0] ));
 dfrtp_2 _24055_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_00992_),
    .RESET_B(net1225),
    .Q(\digitop_pav2.pie_inst.fsm.state[1] ));
 dfrtp_4 _24056_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00993_),
    .RESET_B(net1199),
    .Q(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[0] ));
 dfrtp_4 _24057_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00994_),
    .RESET_B(net1199),
    .Q(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[1] ));
 dfrtp_4 _24058_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00995_),
    .RESET_B(net1199),
    .Q(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[2] ));
 dfrtp_2 _24059_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00996_),
    .RESET_B(net1199),
    .Q(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[3] ));
 dfrtp_2 _24060_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00997_),
    .RESET_B(net1199),
    .Q(\digitop_pav2.invent_inst.invent_tx_pav2.tx_ctr[4] ));
 dfrtp_1 _24061_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00998_),
    .RESET_B(_00236_),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdctr.par4_en_ff ));
 dfrtp_2 _24062_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_00999_),
    .RESET_B(net1454),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.timeout_en_t1 ));
 dfrtp_1 _24063_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01000_),
    .RESET_B(net1447),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmd_abort_b ));
 dfrtp_4 _24064_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01001_),
    .RESET_B(net1447),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.mode ));
 dfrtp_1 _24065_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01002_),
    .RESET_B(net1450),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.piex_dt_rx_done ));
 dfrtp_1 _24066_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(\digitop_pav2.proc_ctrl_inst.cmdfsm.n_crc_eval ),
    .RESET_B(net1439),
    .Q(\digitop_pav2.crc_eval ));
 dfrtp_1 _24067_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01003_),
    .RESET_B(net1447),
    .Q(\digitop_pav2.access_inst.access_ctrl0.f_access_i ));
 dfrtp_1 _24068_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(\digitop_pav2.proc_ctrl_inst.cmdfsm.n_rn_rst_b ),
    .RESET_B(net1441),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.rn_rst_b ));
 dfrtp_1 _24069_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(\digitop_pav2.proc_ctrl_inst.cmdfsm.n_rn_en ),
    .RESET_B(net1447),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.rn_en ));
 dfrtp_1 _24070_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01004_),
    .RESET_B(net1450),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[0] ));
 dfrtp_1 _24071_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01005_),
    .RESET_B(net1450),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[1] ));
 dfrtp_1 _24072_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01006_),
    .RESET_B(net1451),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[2] ));
 dfstp_1 _24073_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01007_),
    .SET_B(net1451),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[3] ));
 dfrtp_1 _24074_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01008_),
    .RESET_B(net1451),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[4] ));
 dfrtp_1 _24075_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01009_),
    .RESET_B(net1450),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[5] ));
 dfstp_1 _24076_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01010_),
    .SET_B(net1450),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[6] ));
 dfrtp_1 _24077_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01011_),
    .RESET_B(net1451),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[7] ));
 dfrtp_1 _24078_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01012_),
    .RESET_B(net1455),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[8] ));
 dfrtp_1 _24079_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01013_),
    .RESET_B(net1451),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.trcal[9] ));
 dfstp_1 _24080_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01014_),
    .SET_B(net1450),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_trext ));
 dfrtp_1 _24081_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01015_),
    .RESET_B(net1450),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_m[0] ));
 dfrtp_1 _24082_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01016_),
    .RESET_B(net1450),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_m[1] ));
 dfrtp_1 _24083_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01017_),
    .RESET_B(net1451),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.query_dr ));
 dfrtp_1 _24084_ (.CLK(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate1.ck_out ),
    .D(_01018_),
    .RESET_B(net1439),
    .Q(\digitop_pav2.fg_tc ));
 dfrtp_1 _24085_ (.CLK(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate1.ck_out ),
    .D(_01019_),
    .RESET_B(net1439),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_cgen.fg_tc_rx_i ));
 dfrtp_2 _24086_ (.CLK(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate1.ck_out ),
    .D(_01020_),
    .RESET_B(net1439),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_cgen.en_g_sec_i ));
 dfrtp_1 _24087_ (.CLK(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate2.ck_out ),
    .D(_01021_),
    .RESET_B(net1448),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.ebv_rst_b ));
 dfrtp_1 _24088_ (.CLK(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate2.ck_out ),
    .D(_01022_),
    .RESET_B(net1448),
    .Q(\digitop_pav2.proc_ctrl_inst.cmdfsm.ebv_en ));
 dfrtp_1 _24089_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(\digitop_pav2.proc_ctrl_inst.profsm.n_blf_abort ),
    .RESET_B(net1450),
    .Q(\digitop_pav2.proc_ctrl_inst.blf_abort ));
 dfrtp_1 _24090_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01023_),
    .RESET_B(net1243),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.dif ));
 dfrtp_1 _24091_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01024_),
    .RESET_B(net1452),
    .Q(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[0] ));
 dfrtp_2 _24092_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01025_),
    .RESET_B(net1447),
    .Q(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[1] ));
 dfrtp_4 _24093_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01026_),
    .RESET_B(net1447),
    .Q(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[2] ));
 dfrtp_1 _24094_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01027_),
    .RESET_B(net1447),
    .Q(\digitop_pav2.proc_ctrl_inst.profsm.skip_abort ));
 dfrtp_2 _24095_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01028_),
    .RESET_B(net1447),
    .Q(\digitop_pav2.proc_ctrl_inst.profsm.r1_ff ));
 dfxtp_1 _24096_ (.CLK(_00237_),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.neg_i[1] ));
 dfxtp_1 _24097_ (.CLK(_00238_),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.neg_i[2] ));
 dfxtp_1 _24098_ (.CLK(_00239_),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.neg_i[3] ));
 dfxtp_1 _24099_ (.CLK(_00240_),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.neg_i[4] ));
 dfxtp_1 _24100_ (.CLK(_00241_),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.neg_i[5] ));
 dfxtp_1 _24101_ (.CLK(_00242_),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.neg_i[6] ));
 dfxtp_1 _24102_ (.CLK(_00243_),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.neg_i[7] ));
 dfxtp_1 _24103_ (.CLK(_00244_),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.neg_i[8] ));
 dfxtp_1 _24104_ (.CLK(_00245_),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.neg_i[9] ));
 dfstp_1 _24105_ (.CLK(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.Y ),
    .D(_00140_),
    .SET_B(\digitop_pav2.pie_inst.ctr.en_ctr_after_buf ),
    .Q(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.A ));
 dfstp_1 _24106_ (.CLK(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.Y ),
    .D(_00138_),
    .SET_B(\digitop_pav2.pie_inst.ctr.en_ctr_after_buf ),
    .Q(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.A ));
 dfstp_1 _24107_ (.CLK(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.Y ),
    .D(_00141_),
    .SET_B(\digitop_pav2.pie_inst.ctr.en_ctr_after_buf ),
    .Q(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.A ));
 dfstp_1 _24108_ (.CLK(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.Y ),
    .D(_00137_),
    .SET_B(\digitop_pav2.pie_inst.ctr.en_ctr_after_buf ),
    .Q(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.A ));
 dfstp_1 _24109_ (.CLK(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.Y ),
    .D(_00142_),
    .SET_B(\digitop_pav2.pie_inst.ctr.en_ctr_after_buf ),
    .Q(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.A ));
 dfstp_1 _24110_ (.CLK(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.Y ),
    .D(_00143_),
    .SET_B(\digitop_pav2.pie_inst.ctr.en_ctr_after_buf ),
    .Q(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.A ));
 dfstp_1 _24111_ (.CLK(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.Y ),
    .D(_00136_),
    .SET_B(\digitop_pav2.pie_inst.ctr.en_ctr_after_buf ),
    .Q(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.A ));
 dfstp_1 _24112_ (.CLK(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.Y ),
    .D(_00139_),
    .SET_B(\digitop_pav2.pie_inst.ctr.en_ctr_after_buf ),
    .Q(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.A ));
 dfstp_1 _24113_ (.CLK(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.Y ),
    .D(_00135_),
    .SET_B(\digitop_pav2.pie_inst.ctr.en_ctr_after_buf ),
    .Q(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.A ));
 dfstp_1 _24114_ (.CLK(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.Y ),
    .D(net1582),
    .SET_B(\digitop_pav2.pie_inst.ctr.en_ctr_after_buf ),
    .Q(\digitop_pav2.pie_inst.ctr.ovf_b ));
 dfstp_1 _24115_ (.CLK(\digitop_pav2.clkx_piex_clk ),
    .D(_00134_),
    .SET_B(\digitop_pav2.pie_inst.ctr.en_ctr_after_buf ),
    .Q(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.A ));
 dfrtp_1 _24116_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(\digitop_pav2.pie_inst.fsm.n_data_en ),
    .RESET_B(net1225),
    .Q(\digitop_pav2.crc_inst.dt_rx_en_i ));
 dfrtp_1 _24117_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01029_),
    .RESET_B(net1225),
    .Q(\digitop_pav2.pie_inst.delend_o ));
 dfrtp_4 _24118_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01030_),
    .RESET_B(net1454),
    .Q(\digitop_pav2.memctrl_inst.extra_dt_i[12] ));
 dfrtp_4 _24119_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01031_),
    .RESET_B(net1454),
    .Q(\digitop_pav2.memctrl_inst.extra_dt_i[13] ));
 dfrtp_4 _24120_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01032_),
    .RESET_B(net1454),
    .Q(\digitop_pav2.memctrl_inst.extra_dt_i[14] ));
 dfrtp_4 _24121_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01033_),
    .RESET_B(net1454),
    .Q(\digitop_pav2.memctrl_inst.extra_dt_i[15] ));
 dfrtp_1 _24122_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01034_),
    .RESET_B(net1454),
    .Q(\digitop_pav2.pie_inst.fsm.trcal[4] ));
 dfrtp_1 _24123_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01035_),
    .RESET_B(net1454),
    .Q(\digitop_pav2.pie_inst.fsm.trcal[5] ));
 dfrtp_1 _24124_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01036_),
    .RESET_B(net1455),
    .Q(\digitop_pav2.pie_inst.fsm.trcal[6] ));
 dfrtp_1 _24125_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01037_),
    .RESET_B(net1454),
    .Q(\digitop_pav2.pie_inst.fsm.trcal[7] ));
 dfrtp_1 _24126_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01038_),
    .RESET_B(net1454),
    .Q(\digitop_pav2.pie_inst.fsm.trcal[8] ));
 dfrtp_1 _24127_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01039_),
    .RESET_B(net1454),
    .Q(\digitop_pav2.pie_inst.fsm.trcal[9] ));
 dfxtp_1 _24128_ (.CLK(\digitop_pav2.pie_inst.fsm.past_clk_i ),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.dif_pos_fix[0] ));
 dfxtp_1 _24129_ (.CLK(\digitop_pav2.pie_inst.fsm.past_clk_i ),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.past_ctr[1] ));
 dfxtp_1 _24130_ (.CLK(\digitop_pav2.pie_inst.fsm.past_clk_i ),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.past_ctr[2] ));
 dfxtp_1 _24131_ (.CLK(\digitop_pav2.pie_inst.fsm.past_clk_i ),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.past_ctr[3] ));
 dfxtp_2 _24132_ (.CLK(\digitop_pav2.pie_inst.fsm.past_clk_i ),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.past_ctr[4] ));
 dfxtp_1 _24133_ (.CLK(\digitop_pav2.pie_inst.fsm.past_clk_i ),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.past_ctr[5] ));
 dfxtp_1 _24134_ (.CLK(\digitop_pav2.pie_inst.fsm.past_clk_i ),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.past_ctr[6] ));
 dfxtp_1 _24135_ (.CLK(\digitop_pav2.pie_inst.fsm.past_clk_i ),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.past_ctr[7] ));
 dfxtp_1 _24136_ (.CLK(\digitop_pav2.pie_inst.fsm.past_clk_i ),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.past_ctr[8] ));
 dfxtp_2 _24137_ (.CLK(\digitop_pav2.pie_inst.fsm.past_clk_i ),
    .D(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.pie_inst.fsm.past_ctr[9] ));
 dfxtp_1 _24138_ (.CLK(\digitop_pav2.pie_inst.fsm.past_clk_i ),
    .D(\digitop_pav2.pie_inst.ctr.ovf_b ),
    .Q(\digitop_pav2.pie_inst.fsm.past_ovf_b ));
 dfstp_1 _24139_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01040_),
    .SET_B(net1420),
    .Q(\digitop_pav2.memctrl_inst.addr_to_reram[0] ));
 dfrtp_2 _24140_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01041_),
    .RESET_B(net1420),
    .Q(\digitop_pav2.memctrl_inst.addr_to_reram[1] ));
 dfrtp_4 _24141_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01042_),
    .RESET_B(net1420),
    .Q(\digitop_pav2.memctrl_inst.addr_to_reram[2] ));
 dfstp_2 _24142_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01043_),
    .SET_B(net1422),
    .Q(\digitop_pav2.memctrl_inst.addr_to_reram[3] ));
 dfstp_1 _24143_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01044_),
    .SET_B(net1423),
    .Q(\digitop_pav2.memctrl_inst.addr_to_reram[4] ));
 dfrtp_1 _24144_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01045_),
    .RESET_B(net1455),
    .Q(\digitop_pav2.pie_inst.fsm.comp_delimiter_ff ));
 dfrtp_1 _24145_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01046_),
    .RESET_B(net1455),
    .Q(\digitop_pav2.pie_inst.fsm.comp_delimiter_ff2 ));
 dfrtp_1 _24146_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(\digitop_pav2.pie_inst.fsm.dif_pos_fix[0] ),
    .RESET_B(net1226),
    .Q(\digitop_pav2.pie_inst.fsm.temptari[0] ));
 dfrtp_1 _24147_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(\digitop_pav2.pie_inst.fsm.dif_pos_fix[1] ),
    .RESET_B(net1225),
    .Q(\digitop_pav2.pie_inst.fsm.temptari[1] ));
 dfrtp_1 _24148_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(\digitop_pav2.pie_inst.fsm.dif_pos_fix[2] ),
    .RESET_B(net1226),
    .Q(\digitop_pav2.pie_inst.fsm.temptari[2] ));
 dfrtp_2 _24149_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(\digitop_pav2.pie_inst.fsm.dif_pos_fix[3] ),
    .RESET_B(net1225),
    .Q(\digitop_pav2.pie_inst.fsm.temptari[3] ));
 dfrtp_2 _24150_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(\digitop_pav2.pie_inst.fsm.dif_pos_fix[4] ),
    .RESET_B(net1225),
    .Q(\digitop_pav2.pie_inst.fsm.temptari[4] ));
 dfrtp_1 _24151_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(\digitop_pav2.pie_inst.fsm.dif_pos_fix[5] ),
    .RESET_B(net1226),
    .Q(\digitop_pav2.pie_inst.fsm.temptari[5] ));
 dfrtp_1 _24152_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(\digitop_pav2.pie_inst.fsm.dif_pos_fix[6] ),
    .RESET_B(net1226),
    .Q(\digitop_pav2.pie_inst.fsm.temptari[6] ));
 dfrtp_2 _24153_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(\digitop_pav2.pie_inst.fsm.dif_pos_fix[7] ),
    .RESET_B(net1226),
    .Q(\digitop_pav2.pie_inst.fsm.temptari[7] ));
 dfrtp_1 _24154_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(\digitop_pav2.pie_inst.fsm.dif_pos_fix[8] ),
    .RESET_B(net1226),
    .Q(\digitop_pav2.pie_inst.fsm.temptari[8] ));
 dfrtp_1 _24155_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(\digitop_pav2.pie_inst.fsm.dif_pos_fix[9] ),
    .RESET_B(net1226),
    .Q(\digitop_pav2.pie_inst.fsm.temptari[9] ));
 dfrtp_1 _24156_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01047_),
    .RESET_B(net1428),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[0] ));
 dfrtp_1 _24157_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01048_),
    .RESET_B(net1426),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[1] ));
 dfrtp_1 _24158_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01049_),
    .RESET_B(net1426),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[2] ));
 dfrtp_1 _24159_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01050_),
    .RESET_B(net1428),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[3] ));
 dfrtp_1 _24160_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01051_),
    .RESET_B(net1428),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[4] ));
 dfrtp_1 _24161_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01052_),
    .RESET_B(net1425),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[5] ));
 dfrtp_1 _24162_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01053_),
    .RESET_B(net1429),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[6] ));
 dfrtp_1 _24163_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01054_),
    .RESET_B(net1429),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[7] ));
 dfrtp_1 _24164_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01055_),
    .RESET_B(net1428),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[8] ));
 dfrtp_1 _24165_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01056_),
    .RESET_B(net1425),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[9] ));
 dfrtp_1 _24166_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01057_),
    .RESET_B(net1428),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[10] ));
 dfrtp_1 _24167_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01058_),
    .RESET_B(net1426),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[11] ));
 dfrtp_4 _24168_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01059_),
    .RESET_B(net1428),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[12] ));
 dfrtp_1 _24169_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01060_),
    .RESET_B(net1428),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[13] ));
 dfrtp_1 _24170_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01061_),
    .RESET_B(net1429),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[14] ));
 dfrtp_1 _24171_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01062_),
    .RESET_B(net1429),
    .Q(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[15] ));
 dfstp_1 _24172_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01063_),
    .SET_B(net1420),
    .Q(\digitop_pav2.memctrl_inst.bit_addr[0] ));
 dfstp_1 _24173_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01064_),
    .SET_B(net1420),
    .Q(\digitop_pav2.memctrl_inst.bit_addr[1] ));
 dfstp_1 _24174_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01065_),
    .SET_B(net1419),
    .Q(\digitop_pav2.memctrl_inst.bit_addr[2] ));
 dfstp_1 _24175_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01066_),
    .SET_B(net1419),
    .Q(\digitop_pav2.memctrl_inst.bit_addr[3] ));
 dfstp_1 _24176_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01067_),
    .SET_B(net1416),
    .Q(\digitop_pav2.memctrl_inst.ctr[0] ));
 dfstp_1 _24177_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01068_),
    .SET_B(net1416),
    .Q(\digitop_pav2.memctrl_inst.ctr[1] ));
 dfstp_1 _24178_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01069_),
    .SET_B(net1416),
    .Q(\digitop_pav2.memctrl_inst.ctr[2] ));
 dfstp_1 _24179_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01070_),
    .SET_B(net1416),
    .Q(\digitop_pav2.memctrl_inst.ctr[3] ));
 dfstp_1 _24180_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01071_),
    .SET_B(net1419),
    .Q(\digitop_pav2.memctrl_inst.ctr[4] ));
 dfstp_1 _24181_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01072_),
    .SET_B(net1427),
    .Q(\digitop_pav2.memctrl_inst.ctr[5] ));
 dfstp_1 _24182_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01073_),
    .SET_B(net1425),
    .Q(\digitop_pav2.memctrl_inst.ctr[6] ));
 dfstp_1 _24183_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01074_),
    .SET_B(net1425),
    .Q(\digitop_pav2.memctrl_inst.ctr[7] ));
 dfrtp_1 _24184_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01075_),
    .RESET_B(net1420),
    .Q(\digitop_pav2.func_reg_wr_en ));
 dfrtp_1 _24185_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(\digitop_pav2.memctrl_inst.n_prog ),
    .RESET_B(net1417),
    .Q(\digitop_pav2.func_rr_prog ));
 dfrtp_1 _24186_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(\digitop_pav2.memctrl_inst.n_erase ),
    .RESET_B(net1417),
    .Q(\digitop_pav2.func_rr_erase ));
 dfrtp_1 _24187_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(\digitop_pav2.memctrl_inst.n_read ),
    .RESET_B(net1419),
    .Q(\digitop_pav2.func_rr_read ));
 dfrtp_1 _24188_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(\digitop_pav2.memctrl_inst.n_bit_addr_allow ),
    .RESET_B(net1420),
    .Q(\digitop_pav2.memctrl_inst.busy_ff ));
 dfrtp_1 _24189_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(net1610),
    .RESET_B(net1419),
    .Q(\digitop_pav2.memctrl_inst.reg_wr_ok_ff ));
 dfrtp_1 _24190_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(\digitop_pav2.memctrl_inst.reg_wr_ok_ff ),
    .RESET_B(net1419),
    .Q(\digitop_pav2.memctrl_inst.reg_wr_ok_ff2 ));
 dfrtp_1 _24191_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01076_),
    .RESET_B(net1420),
    .Q(\digitop_pav2.memctrl_inst.bit_addr_allow ));
 dfbbn_1 _24192_ (.CLK_N(_00248_),
    .D(_01077_),
    .RESET_B(_00246_),
    .SET_B(_00247_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.s1_i ),
    .Q_N(_00170_));
 dfbbn_2 _24193_ (.CLK_N(_00251_),
    .D(_01078_),
    .RESET_B(_00249_),
    .SET_B(_00250_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_r_ff_i ),
    .Q_N(_11504_));
 dfrtp_1 _24194_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01079_),
    .RESET_B(net1285),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[0] ));
 dfrtp_1 _24195_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01080_),
    .RESET_B(net1283),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[1] ));
 dfrtp_1 _24196_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01081_),
    .RESET_B(net1285),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[2] ));
 dfrtp_1 _24197_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01082_),
    .RESET_B(net1283),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[3] ));
 dfrtp_1 _24198_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01083_),
    .RESET_B(net1283),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[4] ));
 dfrtp_1 _24199_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01084_),
    .RESET_B(net1283),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[5] ));
 dfrtp_1 _24200_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01085_),
    .RESET_B(net1285),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_en_ff[6] ));
 dfrtp_1 _24201_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01086_),
    .RESET_B(net1453),
    .Q(\digitop_pav2.invent_inst.s1_r_o ));
 dfbbn_2 _24202_ (.CLK_N(_00254_),
    .D(_01087_),
    .RESET_B(_00252_),
    .SET_B(_00253_),
    .Q(\digitop_pav2.invent_inst.sl_s_ff ),
    .Q_N(_11503_));
 dfbbn_2 _24203_ (.CLK_N(_00257_),
    .D(_01088_),
    .RESET_B(_00255_),
    .SET_B(_00256_),
    .Q(\digitop_pav2.invent_inst.sl_r_ff ),
    .Q_N(_11502_));
 dfbbn_2 _24204_ (.CLK_N(_00260_),
    .D(_01089_),
    .RESET_B(_00258_),
    .SET_B(_00259_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_s_ff_i ),
    .Q_N(_11501_));
 dfrtp_1 _24205_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01090_),
    .RESET_B(net1453),
    .Q(\digitop_pav2.invent_inst.s1_s_o ));
 dfbbn_2 _24206_ (.CLK_N(_00263_),
    .D(_01091_),
    .RESET_B(_00261_),
    .SET_B(_00262_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_s_ff_i ),
    .Q_N(_11500_));
 dfbbn_2 _24207_ (.CLK_N(_00266_),
    .D(_01092_),
    .RESET_B(_00264_),
    .SET_B(_00265_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_r_ff_i ),
    .Q_N(_11499_));
 dfxtp_1 _24208_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01093_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[0] ));
 dfxtp_2 _24209_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01094_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[7] ));
 dfrtp_2 _24210_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01095_),
    .RESET_B(net1199),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[0] ));
 dfrtp_1 _24211_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01096_),
    .RESET_B(net1199),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[1] ));
 dfrtp_1 _24212_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01097_),
    .RESET_B(net1199),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[2] ));
 dfrtp_4 _24213_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01098_),
    .RESET_B(net1199),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[3] ));
 dfrtp_2 _24214_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01099_),
    .RESET_B(net1692),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[4] ));
 dfrtp_1 _24215_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01100_),
    .RESET_B(net1446),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.s0_i ));
 dfrtp_4 _24216_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01101_),
    .RESET_B(net1270),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[0] ));
 dfrtp_1 _24217_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01102_),
    .RESET_B(net1270),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[1] ));
 dfrtp_1 _24218_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01103_),
    .RESET_B(net1270),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[2] ));
 dfrtp_1 _24219_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01104_),
    .RESET_B(net1270),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[3] ));
 dfrtp_4 _24220_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01105_),
    .RESET_B(net1270),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[4] ));
 dfrtp_4 _24221_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01106_),
    .RESET_B(net1270),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[5] ));
 dfrtp_4 _24222_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01107_),
    .RESET_B(net1270),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[6] ));
 dfrtp_1 _24223_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01108_),
    .RESET_B(net1270),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[7] ));
 dfrtp_1 _24224_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01109_),
    .RESET_B(net1271),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[8] ));
 dfxtp_1 _24225_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01110_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[0] ));
 dfxtp_1 _24226_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01111_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[1] ));
 dfxtp_1 _24227_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01112_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[2] ));
 dfxtp_1 _24228_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01113_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[3] ));
 dfxtp_1 _24229_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01114_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[4] ));
 dfxtp_1 _24230_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01115_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[5] ));
 dfxtp_1 _24231_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01116_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[6] ));
 dfxtp_1 _24232_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01117_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[7] ));
 dfxtp_1 _24233_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01118_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[8] ));
 dfxtp_1 _24234_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01119_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[9] ));
 dfxtp_1 _24235_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01120_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[10] ));
 dfxtp_1 _24236_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01121_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[11] ));
 dfxtp_1 _24237_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01122_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[12] ));
 dfxtp_1 _24238_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01123_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[13] ));
 dfxtp_1 _24239_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01124_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[14] ));
 dfxtp_1 _24240_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01125_),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.buf1[15] ));
 dfrtp_4 _24241_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01126_),
    .RESET_B(net1269),
    .Q(\digitop_pav2.invent_inst.invent_sel_pav2.mask_mismatch_ff ));
 dfxtp_1 _24242_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01127_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[0] ));
 dfxtp_1 _24243_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01128_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[1] ));
 dfxtp_1 _24244_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01129_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[2] ));
 dfxtp_1 _24245_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01130_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[3] ));
 dfxtp_1 _24246_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01131_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[4] ));
 dfxtp_1 _24247_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01132_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[5] ));
 dfxtp_1 _24248_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01133_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[6] ));
 dfxtp_1 _24249_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01134_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[7] ));
 dfxtp_1 _24250_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01135_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[8] ));
 dfxtp_1 _24251_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01136_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[9] ));
 dfxtp_1 _24252_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01137_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[10] ));
 dfxtp_1 _24253_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01138_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[11] ));
 dfxtp_1 _24254_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01139_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[12] ));
 dfxtp_1 _24255_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01140_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[13] ));
 dfxtp_1 _24256_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01141_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.slot_ctr[14] ));
 dfstp_1 _24257_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00054_),
    .SET_B(_00267_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[0] ));
 dfrtp_1 _24258_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00058_),
    .RESET_B(net1679),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[1] ));
 dfrtp_1 _24259_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00059_),
    .RESET_B(_00269_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[2] ));
 dfrtp_4 _24260_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00060_),
    .RESET_B(net1673),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[4] ));
 dfrtp_4 _24261_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00061_),
    .RESET_B(net1682),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[6] ));
 dfrtp_1 _24262_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00062_),
    .RESET_B(_00272_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[7] ));
 dfrtp_4 _24263_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00063_),
    .RESET_B(_00273_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.flags_en_o ));
 dfrtp_1 _24264_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00055_),
    .RESET_B(_00274_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.r_invent2_o ));
 dfrtp_2 _24265_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00056_),
    .RESET_B(net1670),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[11] ));
 dfrtp_1 _24266_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_00057_),
    .RESET_B(_00276_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.r_invent3_o ));
 dfxtp_1 _24267_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01142_),
    .Q(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer3_o[7] ));
 dfxtp_1 _24268_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01143_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.query_inversion ));
 dfxtp_2 _24269_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01144_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[0] ));
 dfxtp_1 _24270_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01145_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[1] ));
 dfxtp_1 _24271_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01146_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[2] ));
 dfxtp_2 _24272_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01147_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[3] ));
 dfxtp_1 _24273_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01148_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[0] ));
 dfxtp_1 _24274_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01149_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.prior_session[1] ));
 dfrtp_1 _24275_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(\digitop_pav2.fm0miller_inst.fm0x_ctrl.n_data_valid ),
    .RESET_B(net1283),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.mod_en ));
 dfrtp_1 _24276_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(\digitop_pav2.fm0miller_inst.fm0x_ctrl.n_dt_tx_st ),
    .RESET_B(net1285),
    .Q(\digitop_pav2.fm0miller_inst.dt_tx_st_o ));
 dfstp_1 _24277_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01150_),
    .SET_B(_00277_),
    .Q(\digitop_pav2.crc_inst.crc16_q[0] ));
 dfstp_1 _24278_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01151_),
    .SET_B(_00278_),
    .Q(\digitop_pav2.crc_inst.crc16_q[1] ));
 dfstp_1 _24279_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01152_),
    .SET_B(_00279_),
    .Q(\digitop_pav2.crc_inst.crc16_q[2] ));
 dfstp_1 _24280_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01153_),
    .SET_B(_00280_),
    .Q(\digitop_pav2.crc_inst.crc16_q[3] ));
 dfstp_1 _24281_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01154_),
    .SET_B(_00281_),
    .Q(\digitop_pav2.crc_inst.crc16_q[4] ));
 dfstp_1 _24282_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01155_),
    .SET_B(_00282_),
    .Q(\digitop_pav2.crc_inst.crc16_q[5] ));
 dfstp_1 _24283_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01156_),
    .SET_B(_00283_),
    .Q(\digitop_pav2.crc_inst.crc16_q[6] ));
 dfstp_1 _24284_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01157_),
    .SET_B(_00284_),
    .Q(\digitop_pav2.crc_inst.crc16_q[7] ));
 dfstp_1 _24285_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01158_),
    .SET_B(_00285_),
    .Q(\digitop_pav2.crc_inst.crc16_q[8] ));
 dfstp_1 _24286_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01159_),
    .SET_B(_00286_),
    .Q(\digitop_pav2.crc_inst.crc16_q[9] ));
 dfstp_1 _24287_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01160_),
    .SET_B(_00287_),
    .Q(\digitop_pav2.crc_inst.crc16_q[10] ));
 dfstp_1 _24288_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01161_),
    .SET_B(_00288_),
    .Q(\digitop_pav2.crc_inst.crc16_q[11] ));
 dfstp_1 _24289_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01162_),
    .SET_B(_00289_),
    .Q(\digitop_pav2.crc_inst.crc16_q[12] ));
 dfstp_1 _24290_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01163_),
    .SET_B(_00290_),
    .Q(\digitop_pav2.crc_inst.crc16_q[13] ));
 dfstp_1 _24291_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01164_),
    .SET_B(_00291_),
    .Q(\digitop_pav2.crc_inst.crc16_q[14] ));
 dfstp_1 _24292_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01165_),
    .SET_B(_00292_),
    .Q(\digitop_pav2.crc_inst.crc16_q[15] ));
 dfrtp_1 _24293_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01166_),
    .RESET_B(net1283),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[0] ));
 dfrtp_1 _24294_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01167_),
    .RESET_B(net1283),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[1] ));
 dfrtp_1 _24295_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01168_),
    .RESET_B(net1283),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[2] ));
 dfrtp_2 _24296_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01169_),
    .RESET_B(net1284),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[0] ));
 dfrtp_1 _24297_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01170_),
    .RESET_B(net1285),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[1] ));
 dfrtp_4 _24298_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01171_),
    .RESET_B(net1285),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[2] ));
 dfrtp_4 _24299_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01172_),
    .RESET_B(net1284),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[3] ));
 dfrtp_1 _24300_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01173_),
    .RESET_B(net1284),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[4] ));
 dfrtp_1 _24301_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01174_),
    .RESET_B(net1285),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[0] ));
 dfrtp_1 _24302_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01175_),
    .RESET_B(net1283),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[1] ));
 dfrtp_1 _24303_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01176_),
    .RESET_B(net1283),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.fmctr[2] ));
 dfrtp_1 _24304_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01177_),
    .RESET_B(net1284),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[0] ));
 dfrtp_1 _24305_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01178_),
    .RESET_B(net1284),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[1] ));
 dfrtp_1 _24306_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01179_),
    .RESET_B(net1284),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[2] ));
 dfrtp_1 _24307_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01180_),
    .RESET_B(net1284),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[3] ));
 dfrtp_1 _24308_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01181_),
    .RESET_B(net1284),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[4] ));
 dfrtp_1 _24309_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01182_),
    .RESET_B(net1284),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[5] ));
 dfrtp_1 _24310_ (.CLK(\digitop_pav2.clkx_fm0x_clk ),
    .D(_01183_),
    .RESET_B(net1284),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_ctrl.dt_ff[6] ));
 dfrtp_1 _24311_ (.CLK(_00293_),
    .D(\digitop_pav2.fm0miller_inst.fm0x_ctrl.n_gor ),
    .RESET_B(net192),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[0].fm0miller_pav2_gor_dly.A ));
 dfstp_1 _24312_ (.CLK(_00294_),
    .D(\digitop_pav2.fm0miller_inst.fm0x_ctrl.n_gand ),
    .SET_B(net192),
    .Q(\digitop_pav2.fm0miller_inst.fm0x_mask.gand ));
 dfxtp_1 _24313_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01184_),
    .Q(\digitop_pav2.crc_inst.mctrl_data_end_ff ));
 dfrtp_1 _24314_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01185_),
    .RESET_B(_00295_),
    .Q(\digitop_pav2.crc_inst.count[0] ));
 dfrtp_1 _24315_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01186_),
    .RESET_B(_00296_),
    .Q(\digitop_pav2.crc_inst.count[1] ));
 dfrtp_1 _24316_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01187_),
    .RESET_B(_00297_),
    .Q(\digitop_pav2.crc_inst.count[2] ));
 dfrtp_1 _24317_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01188_),
    .RESET_B(_00298_),
    .Q(\digitop_pav2.crc_inst.count[3] ));
 dfstp_1 _24318_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01189_),
    .SET_B(_00299_),
    .Q(\digitop_pav2.crc_inst.crc5_q[0] ));
 dfrtp_1 _24319_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01190_),
    .RESET_B(_00300_),
    .Q(\digitop_pav2.crc_inst.crc5_q[1] ));
 dfrtp_1 _24320_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01191_),
    .RESET_B(_00301_),
    .Q(\digitop_pav2.crc_inst.crc5_q[2] ));
 dfstp_1 _24321_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01192_),
    .SET_B(_00302_),
    .Q(\digitop_pav2.crc_inst.crc5_q[3] ));
 dfrtp_1 _24322_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01193_),
    .RESET_B(_00303_),
    .Q(\digitop_pav2.crc_inst.crc5_q[4] ));
 dfstp_1 _24323_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01194_),
    .SET_B(net1439),
    .Q(\digitop_pav2.crc_inst.pie_data_en_ff ));
 dfxtp_1 _24324_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01195_),
    .Q(\digitop_pav2.crc_inst.mctrl_data_en_ff ));
 dfstp_1 _24325_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01196_),
    .SET_B(net1418),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[0] ));
 dfrtp_1 _24326_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01197_),
    .RESET_B(net1418),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[1] ));
 dfrtp_1 _24327_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01198_),
    .RESET_B(net1414),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[2] ));
 dfrtp_1 _24328_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01199_),
    .RESET_B(net1414),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[3] ));
 dfrtp_1 _24329_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01200_),
    .RESET_B(net1418),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[4] ));
 dfrtp_1 _24330_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01201_),
    .RESET_B(net1418),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[5] ));
 dfrtp_1 _24331_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01202_),
    .RESET_B(net1414),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[6] ));
 dfrtp_1 _24332_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01203_),
    .RESET_B(net1414),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[7] ));
 dfrtp_1 _24333_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01204_),
    .RESET_B(net1414),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[8] ));
 dfrtp_1 _24334_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01205_),
    .RESET_B(net1414),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.pctr[9] ));
 dfxtp_1 _24335_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01206_),
    .Q(\digitop_pav2.crc_inst.dt_tx_en_aux ));
 dfrtp_1 _24336_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01207_),
    .RESET_B(net1416),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.en_pctr ));
 dfxtp_1 _24337_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01208_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[0] ));
 dfxtp_1 _24338_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01209_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[1] ));
 dfxtp_1 _24339_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01210_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[2] ));
 dfxtp_2 _24340_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01211_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[3] ));
 dfxtp_1 _24341_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01212_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[4] ));
 dfxtp_2 _24342_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01213_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[5] ));
 dfxtp_2 _24343_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01214_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[6] ));
 dfxtp_2 _24344_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01215_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[7] ));
 dfxtp_2 _24345_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01216_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[8] ));
 dfxtp_2 _24346_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01217_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[9] ));
 dfxtp_4 _24347_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01218_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[10] ));
 dfxtp_2 _24348_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01219_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[11] ));
 dfxtp_2 _24349_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01220_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[12] ));
 dfxtp_2 _24350_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01221_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[13] ));
 dfxtp_2 _24351_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01222_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[14] ));
 dfxtp_2 _24352_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01223_),
    .Q(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[15] ));
 dfrtp_2 _24353_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_state[0] ),
    .RESET_B(net1424),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[0] ));
 dfrtp_4 _24354_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_state[1] ),
    .RESET_B(net1424),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[1] ));
 dfrtp_2 _24355_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_state[2] ),
    .RESET_B(net1416),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[2] ));
 dfrtp_1 _24356_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_state[3] ),
    .RESET_B(net1424),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[3] ));
 dfrtp_1 _24357_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_rd_stb ),
    .RESET_B(net1436),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.nvm_calx_rd_stb_o ));
 dfrtp_1 _24358_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_end_stab_clk ),
    .RESET_B(net1415),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.end_stab_clk_i ));
 dfrtp_1 _24359_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_wr_stb ),
    .RESET_B(net1424),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.nvm_calx_wr_stb_o ));
 dfstp_2 _24360_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01224_),
    .SET_B(net1417),
    .Q(\digitop_pav2.cal_inst.calx_mux.dtest_trim_0_i ));
 dfstp_1 _24361_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01225_),
    .SET_B(net1424),
    .Q(\digitop_pav2.cal_inst.calx_mux.dtest_trim_1_i ));
 dfrtp_4 _24362_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(_01226_),
    .RESET_B(net1424),
    .Q(\digitop_pav2.cal_inst.calx_mux.dtest_trim_2_i ));
 dfrtp_2 _24363_ (.CLK(\digitop_pav2.cal_inst.calx_clk_o ),
    .D(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.n_end ),
    .RESET_B(net1415),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.calx_end_o ));
 dfrtp_1 _24364_ (.CLK(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.auxclk_after_buf ),
    .D(_00131_),
    .RESET_B(net1411),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk2 ));
 dfstp_1 _24365_ (.CLK(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk_dftmux.dft_rp_and ),
    .D(net1583),
    .SET_B(net1415),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.stab_clk_dis ));
 dfrtp_1 _24366_ (.CLK(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk2_after_buf ),
    .D(_00132_),
    .RESET_B(net1411),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk4 ));
 dfrtp_1 _24367_ (.CLK(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.ck_in ),
    .D(net1503),
    .RESET_B(net1415),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.rp_ff[0] ));
 dfrtp_4 _24368_ (.CLK(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.ck_in ),
    .D(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.rp_ff[0] ),
    .RESET_B(net1415),
    .Q(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.ref_pulse_sync_o ));
 dfrtp_4 _24369_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_replay_o ),
    .RESET_B(net1433),
    .Q(\digitop_pav2.boot_inst.r_boot_ff ));
 dfrtp_1 _24370_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01227_),
    .RESET_B(net1445),
    .Q(\digitop_pav2.boot_inst.boot_ctrl0.prev_busy ));
 dfxtp_2 _24371_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01228_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[0] ));
 dfxtp_2 _24372_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01229_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[1] ));
 dfxtp_1 _24373_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01230_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[2] ));
 dfxtp_2 _24374_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01231_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[3] ));
 dfxtp_2 _24375_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01232_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[4] ));
 dfxtp_1 _24376_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01233_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[5] ));
 dfxtp_1 _24377_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01234_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[6] ));
 dfxtp_1 _24378_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01235_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[7] ));
 dfxtp_2 _24379_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01236_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[8] ));
 dfxtp_1 _24380_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01237_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[9] ));
 dfxtp_1 _24381_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01238_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[10] ));
 dfxtp_2 _24382_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01239_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[11] ));
 dfxtp_2 _24383_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01240_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[12] ));
 dfxtp_2 _24384_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01241_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[13] ));
 dfxtp_1 _24385_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01242_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[14] ));
 dfxtp_1 _24386_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01243_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key0_r[15] ));
 dfstp_1 _24387_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01244_),
    .SET_B(net1431),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_stage[0] ));
 dfstp_1 _24388_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01245_),
    .SET_B(net1431),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_stage[1] ));
 dfrtp_2 _24389_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01246_),
    .RESET_B(net1433),
    .Q(\digitop_pav2.boot_inst.boot_ctrl0.act_state_i ));
 dfrtp_2 _24390_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01247_),
    .RESET_B(net1413),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[0] ));
 dfrtp_4 _24391_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01248_),
    .RESET_B(net1413),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[1] ));
 dfrtp_4 _24392_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01249_),
    .RESET_B(net1413),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[2] ));
 dfrtp_4 _24393_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01250_),
    .RESET_B(net1425),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[3] ));
 dfrtp_2 _24394_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01251_),
    .RESET_B(net1425),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[4] ));
 dfrtp_4 _24395_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01252_),
    .RESET_B(net1424),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[5] ));
 dfrtp_2 _24396_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01253_),
    .RESET_B(net1427),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[6] ));
 dfrtp_4 _24397_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01254_),
    .RESET_B(net1424),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[7] ));
 dfrtp_4 _24398_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01255_),
    .RESET_B(net1425),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[8] ));
 dfrtp_4 _24399_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01256_),
    .RESET_B(net1424),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[9] ));
 dfrtp_4 _24400_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01257_),
    .RESET_B(net1413),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[10] ));
 dfrtp_4 _24401_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01258_),
    .RESET_B(net1427),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[11] ));
 dfrtp_1 _24402_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01259_),
    .RESET_B(net1436),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_fg[12] ));
 dfrtp_4 _24403_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01260_),
    .RESET_B(net1424),
    .Q(\digitop_pav2.access_inst.access_check0.fg_i[13] ));
 dfrtp_4 _24404_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01261_),
    .RESET_B(net1433),
    .Q(\digitop_pav2.access_inst.access_check0.permalock_tid_i ));
 dfrtp_2 _24405_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01262_),
    .RESET_B(net1433),
    .Q(\digitop_pav2.boot_inst.boot_ctrl0.proc_boot_end_i ));
 dfstp_1 _24406_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01263_),
    .SET_B(net1435),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[16] ));
 dfrtp_1 _24407_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01264_),
    .RESET_B(net1435),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[17] ));
 dfrtp_1 _24408_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01265_),
    .RESET_B(net1432),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[18] ));
 dfrtp_1 _24409_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01266_),
    .RESET_B(net1434),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[19] ));
 dfrtp_1 _24410_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01267_),
    .RESET_B(net1434),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[20] ));
 dfrtp_1 _24411_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01268_),
    .RESET_B(net1431),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[21] ));
 dfrtp_1 _24412_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01269_),
    .RESET_B(net1434),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[22] ));
 dfstp_1 _24413_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01270_),
    .SET_B(net1434),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[23] ));
 dfrtp_1 _24414_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01271_),
    .RESET_B(net1435),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[24] ));
 dfstp_1 _24415_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01272_),
    .SET_B(net1435),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[25] ));
 dfrtp_1 _24416_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01273_),
    .RESET_B(net1434),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[26] ));
 dfrtp_1 _24417_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01274_),
    .RESET_B(net1434),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[27] ));
 dfrtp_1 _24418_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01275_),
    .RESET_B(net1435),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[28] ));
 dfstp_1 _24419_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01276_),
    .SET_B(net1435),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[29] ));
 dfstp_1 _24420_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01277_),
    .SET_B(net1435),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[30] ));
 dfstp_1 _24421_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01278_),
    .SET_B(net1445),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_mask[31] ));
 dfrtp_1 _24422_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01279_),
    .RESET_B(net1432),
    .Q(\digitop_pav2.boot_inst.boot_ctrl0.replay ));
 dfrtp_1 _24423_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01280_),
    .RESET_B(net1433),
    .Q(\digitop_pav2.boot_inst.boot_proc0.proc_boot_sync ));
 dfrtp_1 _24424_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_01281_),
    .RESET_B(net1433),
    .Q(\digitop_pav2.boot_inst.boot_ctrl0.proc_crc_end_i ));
 dfxtp_1 _24425_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01282_),
    .Q(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_0.A ));
 dfxtp_1 _24426_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01283_),
    .Q(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_0.A ));
 dfxtp_2 _24427_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01284_),
    .Q(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[0] ));
 dfxtp_2 _24428_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01285_),
    .Q(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[1] ));
 dfxtp_1 _24429_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01286_),
    .Q(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[2] ));
 dfxtp_1 _24430_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01287_),
    .Q(\digitop_pav2.aes128_inst.aes128_round.round_cnt_r[3] ));
 dfstp_1 _24431_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00007_),
    .SET_B(net1445),
    .Q(\digitop_pav2.boot_inst.boot_ctrl0.state[0] ));
 dfrtp_2 _24432_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00051_),
    .RESET_B(net1445),
    .Q(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_crc_en ));
 dfrtp_1 _24433_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00052_),
    .RESET_B(net1431),
    .Q(\digitop_pav2.boot_inst.boot_ctrl0.state[2] ));
 dfrtp_1 _24434_ (.CLK(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ),
    .D(_00053_),
    .RESET_B(net1445),
    .Q(\digitop_pav2.boot_inst.boot_ctrl0.state[3] ));
 dfxtp_4 _24435_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01288_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[0] ));
 dfxtp_4 _24436_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01289_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[1] ));
 dfxtp_4 _24437_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01290_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[2] ));
 dfxtp_2 _24438_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01291_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[3] ));
 dfxtp_4 _24439_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01292_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[4] ));
 dfxtp_2 _24440_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01293_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[5] ));
 dfxtp_4 _24441_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01294_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[6] ));
 dfxtp_4 _24442_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01295_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ));
 dfxtp_2 _24443_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01296_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[0] ));
 dfxtp_2 _24444_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01297_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[1] ));
 dfxtp_1 _24445_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01298_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[2] ));
 dfxtp_2 _24446_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01299_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[3] ));
 dfxtp_2 _24447_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01300_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[4] ));
 dfxtp_2 _24448_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01301_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[5] ));
 dfxtp_2 _24449_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01302_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[6] ));
 dfxtp_1 _24450_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01303_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[7] ));
 dfxtp_2 _24451_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01304_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[8] ));
 dfxtp_2 _24452_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01305_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[9] ));
 dfxtp_2 _24453_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01306_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[10] ));
 dfxtp_2 _24454_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01307_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[11] ));
 dfxtp_2 _24455_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01308_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[12] ));
 dfxtp_2 _24456_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01309_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[13] ));
 dfxtp_2 _24457_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01310_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[14] ));
 dfxtp_2 _24458_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01311_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key4_r[15] ));
 dfxtp_2 _24459_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01312_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[0] ));
 dfxtp_2 _24460_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01313_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[1] ));
 dfxtp_2 _24461_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01314_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[2] ));
 dfxtp_2 _24462_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01315_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[3] ));
 dfxtp_2 _24463_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01316_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[4] ));
 dfxtp_2 _24464_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01317_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[5] ));
 dfxtp_1 _24465_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01318_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[6] ));
 dfxtp_1 _24466_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01319_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[7] ));
 dfxtp_1 _24467_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01320_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[8] ));
 dfxtp_1 _24468_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01321_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[9] ));
 dfxtp_1 _24469_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01322_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[10] ));
 dfxtp_1 _24470_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01323_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[11] ));
 dfxtp_1 _24471_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01324_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[12] ));
 dfxtp_1 _24472_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01325_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[13] ));
 dfxtp_1 _24473_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01326_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[14] ));
 dfxtp_1 _24474_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01327_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key3_r[15] ));
 dfxtp_1 _24475_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01328_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[0] ));
 dfxtp_1 _24476_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01329_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[1] ));
 dfxtp_1 _24477_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01330_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[2] ));
 dfxtp_1 _24478_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01331_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[3] ));
 dfxtp_1 _24479_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01332_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[4] ));
 dfxtp_1 _24480_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01333_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[5] ));
 dfxtp_1 _24481_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01334_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[6] ));
 dfxtp_1 _24482_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01335_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[7] ));
 dfxtp_1 _24483_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01336_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[8] ));
 dfxtp_1 _24484_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01337_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[9] ));
 dfxtp_1 _24485_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01338_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[10] ));
 dfxtp_1 _24486_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01339_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[11] ));
 dfxtp_1 _24487_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01340_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[12] ));
 dfxtp_1 _24488_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01341_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[13] ));
 dfxtp_1 _24489_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01342_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[14] ));
 dfxtp_1 _24490_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01343_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key2_r[15] ));
 dfxtp_2 _24491_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01344_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[0] ));
 dfxtp_1 _24492_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01345_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[1] ));
 dfxtp_1 _24493_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01346_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[2] ));
 dfxtp_2 _24494_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01347_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[3] ));
 dfxtp_1 _24495_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01348_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[4] ));
 dfxtp_2 _24496_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01349_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[5] ));
 dfxtp_1 _24497_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01350_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[6] ));
 dfxtp_1 _24498_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01351_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[7] ));
 dfxtp_1 _24499_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01352_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[8] ));
 dfxtp_1 _24500_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01353_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[9] ));
 dfxtp_1 _24501_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01354_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[10] ));
 dfxtp_1 _24502_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01355_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[11] ));
 dfxtp_1 _24503_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01356_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[12] ));
 dfxtp_1 _24504_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01357_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[13] ));
 dfxtp_1 _24505_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01358_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[14] ));
 dfxtp_1 _24506_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01359_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key1_r[15] ));
 dfxtp_2 _24507_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01360_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[0] ));
 dfxtp_2 _24508_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01361_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[1] ));
 dfxtp_2 _24509_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01362_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[2] ));
 dfxtp_2 _24510_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01363_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[3] ));
 dfxtp_2 _24511_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01364_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[4] ));
 dfxtp_1 _24512_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01365_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[5] ));
 dfxtp_1 _24513_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01366_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[6] ));
 dfxtp_2 _24514_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01367_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[7] ));
 dfxtp_1 _24515_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01368_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[8] ));
 dfxtp_1 _24516_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01369_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[9] ));
 dfxtp_1 _24517_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01370_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[10] ));
 dfxtp_1 _24518_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01371_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[11] ));
 dfxtp_2 _24519_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01372_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[12] ));
 dfxtp_1 _24520_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01373_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[13] ));
 dfxtp_1 _24521_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01374_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[14] ));
 dfxtp_1 _24522_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01375_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key7_r[15] ));
 dfxtp_2 _24523_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01376_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[0] ));
 dfxtp_1 _24524_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01377_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[1] ));
 dfxtp_2 _24525_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01378_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[2] ));
 dfxtp_1 _24526_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01379_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[3] ));
 dfxtp_1 _24527_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01380_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[4] ));
 dfxtp_1 _24528_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01381_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[5] ));
 dfxtp_1 _24529_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01382_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[6] ));
 dfxtp_1 _24530_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01383_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[7] ));
 dfxtp_1 _24531_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01384_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[8] ));
 dfxtp_1 _24532_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01385_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[9] ));
 dfxtp_1 _24533_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01386_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[10] ));
 dfxtp_2 _24534_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01387_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[11] ));
 dfxtp_1 _24535_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01388_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[12] ));
 dfxtp_1 _24536_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01389_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[13] ));
 dfxtp_1 _24537_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01390_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[14] ));
 dfxtp_1 _24538_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01391_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key6_r[15] ));
 dfxtp_2 _24539_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01392_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[0] ));
 dfxtp_2 _24540_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01393_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[1] ));
 dfxtp_1 _24541_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01394_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[2] ));
 dfxtp_1 _24542_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01395_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[3] ));
 dfxtp_2 _24543_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01396_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[4] ));
 dfxtp_1 _24544_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01397_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[5] ));
 dfxtp_2 _24545_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01398_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[6] ));
 dfxtp_1 _24546_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01399_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[7] ));
 dfxtp_1 _24547_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01400_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[8] ));
 dfxtp_2 _24548_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01401_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[9] ));
 dfxtp_1 _24549_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01402_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[10] ));
 dfxtp_1 _24550_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01403_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[11] ));
 dfxtp_1 _24551_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01404_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[12] ));
 dfxtp_1 _24552_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01405_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[13] ));
 dfxtp_1 _24553_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01406_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[14] ));
 dfxtp_1 _24554_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01407_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.key5_r[15] ));
 dfxtp_4 _24555_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01408_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[0] ));
 dfxtp_4 _24556_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01409_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[1] ));
 dfxtp_4 _24557_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01410_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ));
 dfxtp_2 _24558_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01411_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[3] ));
 dfxtp_2 _24559_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01412_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[4] ));
 dfxtp_2 _24560_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01413_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[5] ));
 dfxtp_2 _24561_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01414_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[6] ));
 dfxtp_4 _24562_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01415_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ));
 dfxtp_2 _24563_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01416_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[8] ));
 dfxtp_2 _24564_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01417_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[9] ));
 dfxtp_4 _24565_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01418_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[10] ));
 dfxtp_2 _24566_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01419_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[11] ));
 dfxtp_2 _24567_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01420_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[12] ));
 dfxtp_2 _24568_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01421_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[13] ));
 dfxtp_2 _24569_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01422_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[14] ));
 dfxtp_2 _24570_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01423_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state1_r[15] ));
 dfxtp_4 _24571_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01424_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[8] ));
 dfxtp_4 _24572_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01425_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[9] ));
 dfxtp_4 _24573_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01426_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[10] ));
 dfxtp_2 _24574_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01427_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[11] ));
 dfxtp_4 _24575_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01428_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[12] ));
 dfxtp_2 _24576_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01429_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[13] ));
 dfxtp_2 _24577_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01430_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[14] ));
 dfxtp_4 _24578_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01431_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state2_r[15] ));
 dfxtp_2 _24579_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01432_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[8] ));
 dfxtp_2 _24580_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01433_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[9] ));
 dfxtp_4 _24581_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01434_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[10] ));
 dfxtp_2 _24582_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01435_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[11] ));
 dfxtp_2 _24583_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01436_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[12] ));
 dfxtp_2 _24584_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01437_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[13] ));
 dfxtp_2 _24585_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01438_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[14] ));
 dfxtp_2 _24586_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01439_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state3_r[15] ));
 dfxtp_2 _24587_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01440_),
    .Q(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[0] ));
 dfxtp_1 _24588_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01441_),
    .Q(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[1] ));
 dfxtp_2 _24589_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01442_),
    .Q(\digitop_pav2.aes128_inst.aes128_counter.counter_3b_o[2] ));
 dfxtp_2 _24590_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01443_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[8] ));
 dfxtp_1 _24591_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01444_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[9] ));
 dfxtp_4 _24592_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01445_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[10] ));
 dfxtp_2 _24593_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01446_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[11] ));
 dfxtp_2 _24594_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01447_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[12] ));
 dfxtp_2 _24595_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01448_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[13] ));
 dfxtp_4 _24596_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01449_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[14] ));
 dfxtp_2 _24597_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01450_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state7_r[15] ));
 dfxtp_4 _24598_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01451_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[0] ));
 dfxtp_4 _24599_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01452_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[1] ));
 dfxtp_2 _24600_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01453_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[2] ));
 dfxtp_2 _24601_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01454_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[3] ));
 dfxtp_2 _24602_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01455_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[4] ));
 dfxtp_2 _24603_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01456_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[5] ));
 dfxtp_2 _24604_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01457_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[6] ));
 dfxtp_2 _24605_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01458_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state6_r[7] ));
 dfxtp_4 _24606_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01459_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ));
 dfxtp_4 _24607_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01460_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[1] ));
 dfxtp_2 _24608_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01461_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[2] ));
 dfxtp_2 _24609_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01462_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[3] ));
 dfxtp_2 _24610_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01463_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[4] ));
 dfxtp_2 _24611_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01464_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[5] ));
 dfxtp_2 _24612_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01465_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[6] ));
 dfxtp_2 _24613_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_01466_),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ));
 dfrtp_1 _24614_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00130_),
    .RESET_B(net1437),
    .Q(\digitop_pav2.aes128_inst.aes128_regs.aes_exe_o ));
 dfrtp_1 _24615_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00128_),
    .RESET_B(net1444),
    .Q(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_key_o ));
 dfrtp_1 _24616_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00129_),
    .RESET_B(net1437),
    .Q(\digitop_pav2.aes128_inst.aes128_counter.cnt_rnd_en_o ));
 dfrtp_2 _24617_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00126_),
    .RESET_B(net1437),
    .Q(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_2b_o ));
 dfrtp_1 _24618_ (.CLK(\digitop_pav2.aes128_inst.aes128_counter.clk_i ),
    .D(_00127_),
    .RESET_B(net1444),
    .Q(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_3b_o ));
 dfrtp_1 _24619_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01467_),
    .RESET_B(net1265),
    .Q(\digitop_pav2.ack_inst.rcnt_ff[0] ));
 dfrtp_1 _24620_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01468_),
    .RESET_B(net1265),
    .Q(\digitop_pav2.ack_inst.rcnt_ff[1] ));
 dfxtp_1 _24621_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01469_),
    .Q(\digitop_pav2.pie_inst.fsm.pivot[0] ));
 dfxtp_2 _24622_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01470_),
    .Q(\digitop_pav2.pie_inst.fsm.pivot[1] ));
 dfxtp_2 _24623_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01471_),
    .Q(\digitop_pav2.pie_inst.fsm.pivot[2] ));
 dfxtp_1 _24624_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01472_),
    .Q(\digitop_pav2.pie_inst.fsm.pivot[3] ));
 dfxtp_2 _24625_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01473_),
    .Q(\digitop_pav2.pie_inst.fsm.pivot[4] ));
 dfxtp_2 _24626_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01474_),
    .Q(\digitop_pav2.pie_inst.fsm.pivot[5] ));
 dfxtp_1 _24627_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01475_),
    .Q(\digitop_pav2.pie_inst.fsm.pivot[6] ));
 dfxtp_2 _24628_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01476_),
    .Q(\digitop_pav2.pie_inst.fsm.pivot[7] ));
 dfxtp_2 _24629_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01477_),
    .Q(\digitop_pav2.pie_inst.fsm.pivot[8] ));
 dfrtp_4 _24630_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01478_),
    .RESET_B(net1264),
    .Q(\digitop_pav2.ack_inst.cnt_ff[0] ));
 dfrtp_1 _24631_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01479_),
    .RESET_B(net1265),
    .Q(\digitop_pav2.ack_inst.cnt_ff[1] ));
 dfrtp_1 _24632_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01480_),
    .RESET_B(net1264),
    .Q(\digitop_pav2.ack_inst.cnt_ff[2] ));
 dfrtp_1 _24633_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01481_),
    .RESET_B(net1264),
    .Q(\digitop_pav2.ack_inst.cnt_ff[3] ));
 dfxtp_1 _24634_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01482_),
    .Q(\digitop_pav2.access_inst.access_check0.wordptr_i[0] ));
 dfxtp_1 _24635_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01483_),
    .Q(\digitop_pav2.access_inst.access_check0.wordptr_i[1] ));
 dfxtp_1 _24636_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01484_),
    .Q(\digitop_pav2.access_inst.access_check0.wordptr_i[2] ));
 dfxtp_1 _24637_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01485_),
    .Q(\digitop_pav2.access_inst.access_check0.wordptr_i[3] ));
 dfxtp_1 _24638_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01486_),
    .Q(\digitop_pav2.access_inst.access_check0.wordptr_i[4] ));
 dfxtp_1 _24639_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01487_),
    .Q(\digitop_pav2.access_inst.access_check0.wordptr_i[5] ));
 dfxtp_1 _24640_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01488_),
    .Q(\digitop_pav2.access_inst.access_check0.wordptr_i[6] ));
 dfrtp_1 _24641_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01489_),
    .RESET_B(net1266),
    .Q(\digitop_pav2.ack_inst.buffer_ff[0] ));
 dfrtp_1 _24642_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01490_),
    .RESET_B(net1264),
    .Q(\digitop_pav2.ack_inst.buffer_ff[1] ));
 dfrtp_1 _24643_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01491_),
    .RESET_B(net1266),
    .Q(\digitop_pav2.ack_inst.buffer_ff[2] ));
 dfrtp_1 _24644_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01492_),
    .RESET_B(net1264),
    .Q(\digitop_pav2.ack_inst.buffer_ff[3] ));
 dfrtp_1 _24645_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01493_),
    .RESET_B(net1266),
    .Q(\digitop_pav2.ack_inst.buffer_ff[4] ));
 dfrtp_1 _24646_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01494_),
    .RESET_B(net1266),
    .Q(\digitop_pav2.ack_inst.buffer_ff[5] ));
 dfrtp_1 _24647_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01495_),
    .RESET_B(net1266),
    .Q(\digitop_pav2.ack_inst.buffer_ff[6] ));
 dfrtp_1 _24648_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01496_),
    .RESET_B(net1264),
    .Q(\digitop_pav2.ack_inst.buffer_ff[7] ));
 dfrtp_1 _24649_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01497_),
    .RESET_B(net1264),
    .Q(\digitop_pav2.ack_inst.buffer_ff[8] ));
 dfrtp_1 _24650_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01498_),
    .RESET_B(net1264),
    .Q(\digitop_pav2.ack_inst.buffer_ff[9] ));
 dfrtp_1 _24651_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01499_),
    .RESET_B(net1266),
    .Q(\digitop_pav2.ack_inst.buffer_ff[10] ));
 dfstp_1 _24652_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01500_),
    .SET_B(net1267),
    .Q(\digitop_pav2.ack_inst.buffer_ff[11] ));
 dfstp_1 _24653_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01501_),
    .SET_B(net1265),
    .Q(\digitop_pav2.ack_inst.buffer_ff[12] ));
 dfrtp_1 _24654_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01502_),
    .RESET_B(net1265),
    .Q(\digitop_pav2.ack_inst.buffer_ff[13] ));
 dfrtp_1 _24655_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01503_),
    .RESET_B(net1265),
    .Q(\digitop_pav2.ack_inst.buffer_ff[14] ));
 dfrtp_1 _24656_ (.CLK(\digitop_pav2.ack_inst.clk_i ),
    .D(_01504_),
    .RESET_B(net1265),
    .Q(\digitop_pav2.ack_inst.buffer_ff[15] ));
 dfrtp_1 _24657_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01505_),
    .RESET_B(_00304_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt ));
 dfrtp_1 _24658_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01506_),
    .RESET_B(_00305_),
    .Q(\digitop_pav2.access_inst.access_check0.wcnt_check_one ));
 dfrtp_2 _24659_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01507_),
    .RESET_B(\digitop_pav2.access_inst.access_check0.permalock_tid_i ),
    .Q(\digitop_pav2.acc_activate ));
 dfrtp_2 _24660_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01508_),
    .RESET_B(_00306_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.replay_ok ));
 dfrtp_4 _24661_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01509_),
    .RESET_B(_00307_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.replay_nok ));
 dfrtp_1 _24662_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01510_),
    .RESET_B(_00308_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.dt_acc_done ));
 dfrtp_1 _24663_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01511_),
    .RESET_B(_00309_),
    .Q(\digitop_pav2.access_inst.access_check0.lock_error_o ));
 dfrtp_1 _24664_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01512_),
    .RESET_B(_00310_),
    .Q(\digitop_pav2.access_inst.access_check0.wr_check_sync_o ));
 dfrtp_1 _24665_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01513_),
    .RESET_B(_00311_),
    .Q(\digitop_pav2.access_inst.access_check0.mem_sign_check_sync_o ));
 dfrtp_2 _24666_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01514_),
    .RESET_B(_00312_),
    .Q(\digitop_pav2.access_inst.access_check0.ctrl_wcknzero_ck ));
 dfrtp_1 _24667_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01515_),
    .RESET_B(_00313_),
    .Q(\digitop_pav2.access_inst.access_check0.write_error_reg ));
 dfrtp_1 _24668_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01516_),
    .RESET_B(net1322),
    .Q(\digitop_pav2.access_inst.acc_wcknzero_o ));
 dfrtp_1 _24669_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01517_),
    .RESET_B(_00314_),
    .Q(\digitop_pav2.access_inst.access_check0.error_word_cnt_ptr ));
 dfrtp_1 _24670_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01518_),
    .RESET_B(\digitop_pav2.access_inst.access_check0.permalock_tid_i ),
    .Q(\digitop_pav2.access_inst.access_check0.act_lock_st ));
 dfrtp_1 _24671_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01519_),
    .RESET_B(_00315_),
    .Q(\digitop_pav2.access_inst.access_check0.pc_invalid_o ));
 dfrtp_1 _24672_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01520_),
    .RESET_B(_00316_),
    .Q(\digitop_pav2.access_inst.access_check0.pc_lock_check_sync_o ));
 dfrtp_1 _24673_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01521_),
    .RESET_B(_00317_),
    .Q(\digitop_pav2.access_inst.access_check0.wcnt_check_zero ));
 dfrtp_1 _24674_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01522_),
    .RESET_B(_00318_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.wr_key_finish_i ));
 dfrtp_1 _24675_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01523_),
    .RESET_B(_00319_),
    .Q(\digitop_pav2.access_inst.access_proc0.ctrl_rd_bus_res ));
 dfrtp_2 _24676_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01524_),
    .RESET_B(_00320_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.prev_busy ));
 dfrtp_1 _24677_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01525_),
    .RESET_B(_00321_),
    .Q(\digitop_pav2.access_inst.access_proc0.ctrl_rd_bus ));
 dfrtp_1 _24678_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01526_),
    .RESET_B(_00322_),
    .Q(\digitop_pav2.access_inst.access_check0.proc_finish1_i ));
 dfrtp_1 _24679_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01527_),
    .RESET_B(_00323_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.ld_dt_env_finish_i ));
 dfrtp_1 _24680_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01528_),
    .RESET_B(_00324_),
    .Q(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[0] ));
 dfrtp_1 _24681_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01529_),
    .RESET_B(_00325_),
    .Q(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[1] ));
 dfrtp_1 _24682_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01530_),
    .RESET_B(_00326_),
    .Q(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[2] ));
 dfrtp_1 _24683_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01531_),
    .RESET_B(_00327_),
    .Q(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[3] ));
 dfrtp_1 _24684_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01532_),
    .RESET_B(_00328_),
    .Q(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[7] ));
 dfrtp_1 _24685_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01533_),
    .RESET_B(_00329_),
    .Q(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[8] ));
 dfrtp_4 _24686_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01534_),
    .RESET_B(_00330_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.crc_init_i ));
 dfrtp_1 _24687_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01535_),
    .RESET_B(_00331_),
    .Q(\digitop_pav2.access_inst.access_proc0.proc_crc_check[0] ));
 dfrtp_4 _24688_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01536_),
    .RESET_B(_00332_),
    .Q(\digitop_pav2.access_inst.access_proc0.proc_crc_check[1] ));
 dfrtp_1 _24689_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01537_),
    .RESET_B(_00333_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.proc_finish0_i ));
 dfrtp_2 _24690_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01538_),
    .RESET_B(_00334_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.ld_key_env_finish_i ));
 dfrtp_4 _24691_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01539_),
    .RESET_B(_00335_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.tx_proc_rd_stb_i ));
 dfrtp_1 _24692_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01540_),
    .RESET_B(_00336_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.ctrl_circ_buf ));
 dfrtp_2 _24693_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01541_),
    .RESET_B(_00337_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[0] ));
 dfrtp_2 _24694_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01542_),
    .RESET_B(_00338_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[1] ));
 dfrtp_1 _24695_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01543_),
    .RESET_B(_00339_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[2] ));
 dfrtp_1 _24696_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01544_),
    .RESET_B(_00340_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[3] ));
 dfrtp_1 _24697_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01545_),
    .RESET_B(_00341_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.tx_bit_i ));
 dfrtp_2 _24698_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01546_),
    .RESET_B(_00342_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.rx_par0_i ));
 dfrtp_1 _24699_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01547_),
    .RESET_B(_00343_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.rx_par1_i ));
 dfrtp_1 _24700_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01548_),
    .RESET_B(_00344_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.tx_dt_finish_i ));
 dfxtp_1 _24701_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01549_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[0] ));
 dfxtp_1 _24702_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01550_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[1] ));
 dfxtp_1 _24703_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01551_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[2] ));
 dfxtp_1 _24704_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01552_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[3] ));
 dfxtp_1 _24705_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01553_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[4] ));
 dfxtp_2 _24706_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01554_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[5] ));
 dfxtp_2 _24707_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01555_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[6] ));
 dfxtp_2 _24708_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01556_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[7] ));
 dfxtp_2 _24709_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01557_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[8] ));
 dfxtp_2 _24710_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01558_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[9] ));
 dfxtp_2 _24711_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01559_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[10] ));
 dfxtp_2 _24712_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01560_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[11] ));
 dfxtp_2 _24713_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01561_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[12] ));
 dfxtp_2 _24714_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01562_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[13] ));
 dfxtp_2 _24715_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01563_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[14] ));
 dfxtp_2 _24716_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01564_),
    .Q(\digitop_pav2.access_inst.access_proc0.access_crc16_prl0.crc16[15] ));
 dfrtp_1 _24717_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01565_),
    .RESET_B(_00345_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.dt_acc_done_o ));
 dfrtp_1 _24718_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01566_),
    .RESET_B(_00346_),
    .Q(\digitop_pav2.access_inst.access_check0.error_wordcnt_i ));
 dfrtp_1 _24719_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01567_),
    .RESET_B(_00347_),
    .Q(\digitop_pav2.access_inst.access_transceiver0.wcnt_stb_valid ));
 dfxtp_2 _24720_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01568_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[0] ));
 dfxtp_2 _24721_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01569_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[1] ));
 dfxtp_2 _24722_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01570_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[2] ));
 dfxtp_2 _24723_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01571_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[3] ));
 dfxtp_2 _24724_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01572_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[4] ));
 dfxtp_2 _24725_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01573_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[5] ));
 dfxtp_2 _24726_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01574_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[6] ));
 dfxtp_2 _24727_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01575_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[7] ));
 dfxtp_2 _24728_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01576_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[8] ));
 dfxtp_2 _24729_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01577_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[9] ));
 dfxtp_2 _24730_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01578_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[10] ));
 dfxtp_2 _24731_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01579_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[11] ));
 dfxtp_2 _24732_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01580_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[12] ));
 dfxtp_2 _24733_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01581_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[13] ));
 dfxtp_1 _24734_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01582_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[14] ));
 dfxtp_1 _24735_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01583_),
    .Q(\digitop_pav2.access_inst.access_check0.rx_wr_dt_to_nvm_i[15] ));
 dfrtp_1 _24736_ (.CLK(\digitop_pav2.access_inst.access_check0.clk_i ),
    .D(_01584_),
    .RESET_B(_00348_),
    .Q(\digitop_pav2.access_inst.access_ctrl0.proc_rd_finish_i ));
 dfrtp_1 _24737_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01585_),
    .RESET_B(net1426),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[0] ));
 dfrtp_1 _24738_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01586_),
    .RESET_B(net1425),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[1] ));
 dfrtp_1 _24739_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01587_),
    .RESET_B(net1426),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[2] ));
 dfrtp_1 _24740_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01588_),
    .RESET_B(net1428),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[3] ));
 dfrtp_1 _24741_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01589_),
    .RESET_B(net1430),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[4] ));
 dfrtp_1 _24742_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01590_),
    .RESET_B(net1426),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[5] ));
 dfrtp_1 _24743_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01591_),
    .RESET_B(net1430),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[6] ));
 dfrtp_1 _24744_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01592_),
    .RESET_B(net1429),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[7] ));
 dfrtp_1 _24745_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01593_),
    .RESET_B(net1423),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[8] ));
 dfrtp_1 _24746_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01594_),
    .RESET_B(net1419),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[9] ));
 dfrtp_1 _24747_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01595_),
    .RESET_B(net1428),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[10] ));
 dfrtp_1 _24748_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01596_),
    .RESET_B(net1428),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[11] ));
 dfrtp_1 _24749_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01597_),
    .RESET_B(net1430),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[12] ));
 dfrtp_1 _24750_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01598_),
    .RESET_B(net1430),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[13] ));
 dfrtp_1 _24751_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01599_),
    .RESET_B(net1429),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[14] ));
 dfrtp_1 _24752_ (.CLK(\digitop_pav2.clkx_mem_top_clk ),
    .D(_01600_),
    .RESET_B(net1429),
    .Q(\digitop_pav2.memctrl_inst.flops_0x081[15] ));
 dfxtp_1 _24753_ (.CLK(\digitop_pav2.pie_inst.fsm.clk_i ),
    .D(_01601_),
    .Q(\digitop_pav2.crc_inst.dt_rx_i ));
 dfrtp_1 _24754_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01602_),
    .RESET_B(net1687),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[13] ));
 dfrtp_1 _24755_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01603_),
    .RESET_B(net1676),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[9] ));
 dfrtp_1 _24756_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01604_),
    .RESET_B(net1684),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[5] ));
 dfrtp_1 _24757_ (.CLK(\digitop_pav2.clkx_invent_clk ),
    .D(_01605_),
    .RESET_B(_00352_),
    .Q(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[3] ));
 dfrtp_1 _24758_ (.CLK(\digitop_pav2.sync_inst.inst_rstx.osc_clk_gated ),
    .D(_01606_),
    .RESET_B(\digitop_pav2.sync_inst.inst_rstx.sync_rstx_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Q(\digitop_pav2.sync_inst.inst_rstx.gray_counter[0] ));
 dfrtp_1 _24759_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01607_),
    .RESET_B(net973),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[14] ));
 dfrtp_1 _24760_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01608_),
    .RESET_B(net973),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[13] ));
 dfrtp_1 _24761_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01609_),
    .RESET_B(net972),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[12] ));
 dfrtp_1 _24762_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01610_),
    .RESET_B(net972),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[11] ));
 dfrtp_1 _24763_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01611_),
    .RESET_B(net973),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[10] ));
 dfrtp_1 _24764_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01612_),
    .RESET_B(net973),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[9] ));
 dfrtp_1 _24765_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01613_),
    .RESET_B(net972),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[7] ));
 dfrtp_1 _24766_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01614_),
    .RESET_B(net972),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[6] ));
 dfrtp_1 _24767_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01615_),
    .RESET_B(net972),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[5] ));
 dfrtp_1 _24768_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01616_),
    .RESET_B(net972),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[3] ));
 dfrtp_1 _24769_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01617_),
    .RESET_B(net973),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[2] ));
 dfrtp_1 _24770_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01618_),
    .RESET_B(net972),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[1] ));
 dfstp_1 _24771_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01619_),
    .SET_B(net972),
    .Q(\digitop_pav2.proc_ctrl_inst.ebv.state[0] ));
 dfrtp_1 _24772_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01620_),
    .RESET_B(net1242),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[15] ));
 dfrtp_1 _24773_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01621_),
    .RESET_B(net1242),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[14] ));
 dfrtp_1 _24774_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01622_),
    .RESET_B(net1242),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[13] ));
 dfrtp_1 _24775_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01623_),
    .RESET_B(net1243),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[12] ));
 dfrtp_1 _24776_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01624_),
    .RESET_B(net1242),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[11] ));
 dfrtp_1 _24777_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01625_),
    .RESET_B(net1242),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[10] ));
 dfrtp_2 _24778_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01626_),
    .RESET_B(net1243),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[9] ));
 dfrtp_1 _24779_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01627_),
    .RESET_B(net1243),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[8] ));
 dfrtp_1 _24780_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01628_),
    .RESET_B(net1242),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[7] ));
 dfrtp_1 _24781_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01629_),
    .RESET_B(net1242),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[6] ));
 dfrtp_1 _24782_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01630_),
    .RESET_B(net1243),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[5] ));
 dfrtp_1 _24783_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01631_),
    .RESET_B(net1242),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[4] ));
 dfrtp_1 _24784_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01632_),
    .RESET_B(net1242),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[3] ));
 dfrtp_1 _24785_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01633_),
    .RESET_B(net1242),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[2] ));
 dfrtp_4 _24786_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01634_),
    .RESET_B(net1243),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[1] ));
 dfstp_1 _24787_ (.CLK(\digitop_pav2.clkx_cp_clk ),
    .D(_01635_),
    .SET_B(net1243),
    .Q(\digitop_pav2.proc_ctrl_inst.inst_checker.state[0] ));
 dfrtp_1 _24788_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_01636_),
    .RESET_B(net1005),
    .Q(\digitop_pav2.sec_inst.ld_mem.st[3] ));
 dfrtp_4 _24789_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_01637_),
    .RESET_B(net1005),
    .Q(\digitop_pav2.sec_inst.ld_mem.st[2] ));
 dfrtp_1 _24790_ (.CLK(\digitop_pav2.clkx_sec_clk ),
    .D(_01638_),
    .RESET_B(net985),
    .Q(\digitop_pav2.sec_inst.shift_out.st[1] ));
 dfrtp_4 _24791_ (.CLK(tclk_i),
    .D(_01639_),
    .RESET_B(net1402),
    .Q(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.form_type[1] ));
 dfrtp_1 _24792_ (.CLK(clk_i),
    .D(_01640_),
    .RESET_B(net1533),
    .Q(\vmem[511] ));
 dfrtp_1 _24793_ (.CLK(clk_i),
    .D(_01641_),
    .RESET_B(net1545),
    .Q(\vmem[510] ));
 dfrtp_1 _24794_ (.CLK(clk_i),
    .D(_01642_),
    .RESET_B(net1556),
    .Q(\vmem[509] ));
 dfrtp_1 _24795_ (.CLK(clk_i),
    .D(_01643_),
    .RESET_B(net1567),
    .Q(\vmem[508] ));
 dfrtp_1 _24796_ (.CLK(clk_i),
    .D(_01644_),
    .RESET_B(net1537),
    .Q(\vmem[507] ));
 dfrtp_1 _24797_ (.CLK(clk_i),
    .D(_01645_),
    .RESET_B(net1521),
    .Q(\vmem[506] ));
 dfrtp_1 _24798_ (.CLK(clk_i),
    .D(_01646_),
    .RESET_B(net1551),
    .Q(\vmem[505] ));
 dfrtp_1 _24799_ (.CLK(clk_i),
    .D(_01647_),
    .RESET_B(net1512),
    .Q(\vmem[504] ));
 dfrtp_1 _24800_ (.CLK(clk_i),
    .D(_01648_),
    .RESET_B(net1529),
    .Q(\vmem[503] ));
 dfrtp_1 _24801_ (.CLK(clk_i),
    .D(_01649_),
    .RESET_B(net1569),
    .Q(\vmem[502] ));
 dfrtp_1 _24802_ (.CLK(clk_i),
    .D(_01650_),
    .RESET_B(net1518),
    .Q(\vmem[501] ));
 dfrtp_1 _24803_ (.CLK(clk_i),
    .D(_01651_),
    .RESET_B(net1556),
    .Q(\vmem[500] ));
 dfrtp_1 _24804_ (.CLK(clk_i),
    .D(_01652_),
    .RESET_B(net1506),
    .Q(\vmem[499] ));
 dfrtp_1 _24805_ (.CLK(clk_i),
    .D(_01653_),
    .RESET_B(net1565),
    .Q(\vmem[498] ));
 dfrtp_1 _24806_ (.CLK(clk_i),
    .D(_01654_),
    .RESET_B(net1576),
    .Q(\vmem[497] ));
 dfrtp_1 _24807_ (.CLK(clk_i),
    .D(_01655_),
    .RESET_B(net1526),
    .Q(\vmem[496] ));
 dfrtp_1 _24808_ (.CLK(clk_i),
    .D(_01656_),
    .RESET_B(net1531),
    .Q(\vmem[495] ));
 dfrtp_1 _24809_ (.CLK(clk_i),
    .D(_01657_),
    .RESET_B(net1560),
    .Q(\vmem[494] ));
 dfrtp_1 _24810_ (.CLK(clk_i),
    .D(_01658_),
    .RESET_B(net1556),
    .Q(\vmem[493] ));
 dfrtp_1 _24811_ (.CLK(clk_i),
    .D(_01659_),
    .RESET_B(net1567),
    .Q(\vmem[492] ));
 dfrtp_1 _24812_ (.CLK(clk_i),
    .D(_01660_),
    .RESET_B(net1537),
    .Q(\vmem[491] ));
 dfrtp_1 _24813_ (.CLK(clk_i),
    .D(_01661_),
    .RESET_B(net1521),
    .Q(\vmem[490] ));
 dfrtp_1 _24814_ (.CLK(clk_i),
    .D(_01662_),
    .RESET_B(net1551),
    .Q(\vmem[489] ));
 dfrtp_1 _24815_ (.CLK(clk_i),
    .D(_01663_),
    .RESET_B(net1512),
    .Q(\vmem[488] ));
 dfrtp_1 _24816_ (.CLK(clk_i),
    .D(_01664_),
    .RESET_B(net1540),
    .Q(\vmem[487] ));
 dfrtp_1 _24817_ (.CLK(clk_i),
    .D(_01665_),
    .RESET_B(net1569),
    .Q(\vmem[486] ));
 dfrtp_1 _24818_ (.CLK(clk_i),
    .D(_01666_),
    .RESET_B(net1518),
    .Q(\vmem[485] ));
 dfrtp_1 _24819_ (.CLK(clk_i),
    .D(_01667_),
    .RESET_B(net1556),
    .Q(\vmem[484] ));
 dfrtp_1 _24820_ (.CLK(clk_i),
    .D(_01668_),
    .RESET_B(net1506),
    .Q(\vmem[483] ));
 dfrtp_1 _24821_ (.CLK(clk_i),
    .D(_01669_),
    .RESET_B(net1558),
    .Q(\vmem[482] ));
 dfrtp_1 _24822_ (.CLK(clk_i),
    .D(_01670_),
    .RESET_B(net1578),
    .Q(\vmem[481] ));
 dfrtp_1 _24823_ (.CLK(clk_i),
    .D(_01671_),
    .RESET_B(net1526),
    .Q(\vmem[480] ));
 dfrtp_1 _24824_ (.CLK(clk_i),
    .D(_01672_),
    .RESET_B(net1533),
    .Q(\vmem[479] ));
 dfrtp_1 _24825_ (.CLK(clk_i),
    .D(_01673_),
    .RESET_B(net1545),
    .Q(\vmem[478] ));
 dfrtp_1 _24826_ (.CLK(clk_i),
    .D(_01674_),
    .RESET_B(net1541),
    .Q(\vmem[477] ));
 dfrtp_1 _24827_ (.CLK(clk_i),
    .D(_01675_),
    .RESET_B(net1567),
    .Q(\vmem[476] ));
 dfrtp_1 _24828_ (.CLK(clk_i),
    .D(_01676_),
    .RESET_B(net1537),
    .Q(\vmem[475] ));
 dfrtp_1 _24829_ (.CLK(clk_i),
    .D(_01677_),
    .RESET_B(net1524),
    .Q(\vmem[474] ));
 dfrtp_1 _24830_ (.CLK(clk_i),
    .D(_01678_),
    .RESET_B(net1551),
    .Q(\vmem[473] ));
 dfrtp_1 _24831_ (.CLK(clk_i),
    .D(_01679_),
    .RESET_B(net1512),
    .Q(\vmem[472] ));
 dfrtp_1 _24832_ (.CLK(clk_i),
    .D(_01680_),
    .RESET_B(net1524),
    .Q(\vmem[471] ));
 dfrtp_1 _24833_ (.CLK(clk_i),
    .D(_01681_),
    .RESET_B(net1570),
    .Q(\vmem[470] ));
 dfrtp_1 _24834_ (.CLK(clk_i),
    .D(_01682_),
    .RESET_B(net1518),
    .Q(\vmem[469] ));
 dfrtp_1 _24835_ (.CLK(clk_i),
    .D(_01683_),
    .RESET_B(net1560),
    .Q(\vmem[468] ));
 dfrtp_1 _24836_ (.CLK(clk_i),
    .D(_01684_),
    .RESET_B(net1507),
    .Q(\vmem[467] ));
 dfrtp_1 _24837_ (.CLK(clk_i),
    .D(_01685_),
    .RESET_B(net1558),
    .Q(\vmem[466] ));
 dfrtp_1 _24838_ (.CLK(clk_i),
    .D(_01686_),
    .RESET_B(net1555),
    .Q(\vmem[465] ));
 dfrtp_1 _24839_ (.CLK(clk_i),
    .D(_01687_),
    .RESET_B(net1526),
    .Q(\vmem[464] ));
 dfrtp_1 _24840_ (.CLK(clk_i),
    .D(_01688_),
    .RESET_B(net1534),
    .Q(\vmem[463] ));
 dfrtp_1 _24841_ (.CLK(clk_i),
    .D(_01689_),
    .RESET_B(net1545),
    .Q(\vmem[462] ));
 dfrtp_1 _24842_ (.CLK(clk_i),
    .D(_01690_),
    .RESET_B(net1541),
    .Q(\vmem[461] ));
 dfrtp_1 _24843_ (.CLK(clk_i),
    .D(_01691_),
    .RESET_B(net1565),
    .Q(\vmem[460] ));
 dfrtp_1 _24844_ (.CLK(clk_i),
    .D(_01692_),
    .RESET_B(net1538),
    .Q(\vmem[459] ));
 dfrtp_1 _24845_ (.CLK(clk_i),
    .D(_01693_),
    .RESET_B(net1524),
    .Q(\vmem[458] ));
 dfrtp_1 _24846_ (.CLK(clk_i),
    .D(_01694_),
    .RESET_B(net1549),
    .Q(\vmem[457] ));
 dfrtp_1 _24847_ (.CLK(clk_i),
    .D(_01695_),
    .RESET_B(net1512),
    .Q(\vmem[456] ));
 dfrtp_1 _24848_ (.CLK(clk_i),
    .D(_01696_),
    .RESET_B(net1524),
    .Q(\vmem[455] ));
 dfrtp_1 _24849_ (.CLK(clk_i),
    .D(_01697_),
    .RESET_B(net1570),
    .Q(\vmem[454] ));
 dfrtp_1 _24850_ (.CLK(clk_i),
    .D(_01698_),
    .RESET_B(net1518),
    .Q(\vmem[453] ));
 dfrtp_1 _24851_ (.CLK(clk_i),
    .D(_01699_),
    .RESET_B(net1560),
    .Q(\vmem[452] ));
 dfrtp_1 _24852_ (.CLK(clk_i),
    .D(_01700_),
    .RESET_B(net1506),
    .Q(\vmem[451] ));
 dfrtp_1 _24853_ (.CLK(clk_i),
    .D(_01701_),
    .RESET_B(net1565),
    .Q(\vmem[450] ));
 dfrtp_1 _24854_ (.CLK(clk_i),
    .D(_01702_),
    .RESET_B(net1567),
    .Q(\vmem[449] ));
 dfrtp_1 _24855_ (.CLK(clk_i),
    .D(_01703_),
    .RESET_B(net1517),
    .Q(\vmem[448] ));
 dfrtp_1 _24856_ (.CLK(clk_i),
    .D(_01704_),
    .RESET_B(net1534),
    .Q(\vmem[447] ));
 dfrtp_1 _24857_ (.CLK(clk_i),
    .D(_01705_),
    .RESET_B(net1546),
    .Q(\vmem[446] ));
 dfrtp_1 _24858_ (.CLK(clk_i),
    .D(_01706_),
    .RESET_B(net1541),
    .Q(\vmem[445] ));
 dfrtp_1 _24859_ (.CLK(clk_i),
    .D(_01707_),
    .RESET_B(net1566),
    .Q(\vmem[444] ));
 dfrtp_1 _24860_ (.CLK(clk_i),
    .D(_01708_),
    .RESET_B(net1538),
    .Q(\vmem[443] ));
 dfrtp_1 _24861_ (.CLK(clk_i),
    .D(_01709_),
    .RESET_B(net1521),
    .Q(\vmem[442] ));
 dfrtp_1 _24862_ (.CLK(clk_i),
    .D(_01710_),
    .RESET_B(net1551),
    .Q(\vmem[441] ));
 dfrtp_1 _24863_ (.CLK(clk_i),
    .D(_01711_),
    .RESET_B(net1512),
    .Q(\vmem[440] ));
 dfrtp_1 _24864_ (.CLK(clk_i),
    .D(_01712_),
    .RESET_B(net1529),
    .Q(\vmem[439] ));
 dfrtp_1 _24865_ (.CLK(clk_i),
    .D(_01713_),
    .RESET_B(net1570),
    .Q(\vmem[438] ));
 dfrtp_1 _24866_ (.CLK(clk_i),
    .D(_01714_),
    .RESET_B(net1518),
    .Q(\vmem[437] ));
 dfrtp_1 _24867_ (.CLK(clk_i),
    .D(_01715_),
    .RESET_B(net1562),
    .Q(\vmem[436] ));
 dfrtp_1 _24868_ (.CLK(clk_i),
    .D(_01716_),
    .RESET_B(net1507),
    .Q(\vmem[435] ));
 dfrtp_1 _24869_ (.CLK(clk_i),
    .D(_01717_),
    .RESET_B(net1558),
    .Q(\vmem[434] ));
 dfrtp_1 _24870_ (.CLK(clk_i),
    .D(_01718_),
    .RESET_B(net1578),
    .Q(\vmem[433] ));
 dfrtp_1 _24871_ (.CLK(clk_i),
    .D(_01719_),
    .RESET_B(net1526),
    .Q(\vmem[432] ));
 dfrtp_1 _24872_ (.CLK(clk_i),
    .D(_01720_),
    .RESET_B(net1532),
    .Q(\vmem[431] ));
 dfrtp_1 _24873_ (.CLK(clk_i),
    .D(_01721_),
    .RESET_B(net1560),
    .Q(\vmem[430] ));
 dfrtp_1 _24874_ (.CLK(clk_i),
    .D(_01722_),
    .RESET_B(net1541),
    .Q(\vmem[429] ));
 dfrtp_1 _24875_ (.CLK(clk_i),
    .D(_01723_),
    .RESET_B(net1568),
    .Q(\vmem[428] ));
 dfrtp_1 _24876_ (.CLK(clk_i),
    .D(_01724_),
    .RESET_B(net1543),
    .Q(\vmem[427] ));
 dfrtp_1 _24877_ (.CLK(clk_i),
    .D(_01725_),
    .RESET_B(net1521),
    .Q(\vmem[426] ));
 dfrtp_1 _24878_ (.CLK(clk_i),
    .D(_01726_),
    .RESET_B(net1551),
    .Q(\vmem[425] ));
 dfrtp_1 _24879_ (.CLK(clk_i),
    .D(_01727_),
    .RESET_B(net1513),
    .Q(\vmem[424] ));
 dfrtp_1 _24880_ (.CLK(clk_i),
    .D(_01728_),
    .RESET_B(net1540),
    .Q(\vmem[423] ));
 dfrtp_1 _24881_ (.CLK(clk_i),
    .D(_01729_),
    .RESET_B(net1571),
    .Q(\vmem[422] ));
 dfrtp_1 _24882_ (.CLK(clk_i),
    .D(_01730_),
    .RESET_B(net1518),
    .Q(\vmem[421] ));
 dfrtp_1 _24883_ (.CLK(clk_i),
    .D(_01731_),
    .RESET_B(net1562),
    .Q(\vmem[420] ));
 dfrtp_1 _24884_ (.CLK(clk_i),
    .D(_01732_),
    .RESET_B(net1507),
    .Q(\vmem[419] ));
 dfrtp_1 _24885_ (.CLK(clk_i),
    .D(_01733_),
    .RESET_B(net1559),
    .Q(\vmem[418] ));
 dfrtp_1 _24886_ (.CLK(clk_i),
    .D(_01734_),
    .RESET_B(net1578),
    .Q(\vmem[417] ));
 dfrtp_1 _24887_ (.CLK(clk_i),
    .D(_01735_),
    .RESET_B(net1526),
    .Q(\vmem[416] ));
 dfrtp_1 _24888_ (.CLK(clk_i),
    .D(_01736_),
    .RESET_B(net1534),
    .Q(\vmem[415] ));
 dfrtp_1 _24889_ (.CLK(clk_i),
    .D(_01737_),
    .RESET_B(net1546),
    .Q(\vmem[414] ));
 dfrtp_1 _24890_ (.CLK(clk_i),
    .D(_01738_),
    .RESET_B(net1541),
    .Q(\vmem[413] ));
 dfrtp_1 _24891_ (.CLK(clk_i),
    .D(_01739_),
    .RESET_B(net1566),
    .Q(\vmem[412] ));
 dfrtp_1 _24892_ (.CLK(clk_i),
    .D(_01740_),
    .RESET_B(net1538),
    .Q(\vmem[411] ));
 dfrtp_1 _24893_ (.CLK(clk_i),
    .D(_01741_),
    .RESET_B(net1522),
    .Q(\vmem[410] ));
 dfrtp_1 _24894_ (.CLK(clk_i),
    .D(_01742_),
    .RESET_B(net1551),
    .Q(\vmem[409] ));
 dfrtp_1 _24895_ (.CLK(clk_i),
    .D(_01743_),
    .RESET_B(net1511),
    .Q(\vmem[408] ));
 dfrtp_1 _24896_ (.CLK(clk_i),
    .D(_01744_),
    .RESET_B(net1533),
    .Q(\vmem[407] ));
 dfrtp_1 _24897_ (.CLK(clk_i),
    .D(_01745_),
    .RESET_B(net1570),
    .Q(\vmem[406] ));
 dfrtp_1 _24898_ (.CLK(clk_i),
    .D(_01746_),
    .RESET_B(net1518),
    .Q(\vmem[405] ));
 dfrtp_1 _24899_ (.CLK(clk_i),
    .D(_01747_),
    .RESET_B(net1560),
    .Q(\vmem[404] ));
 dfrtp_1 _24900_ (.CLK(clk_i),
    .D(_01748_),
    .RESET_B(net1507),
    .Q(\vmem[403] ));
 dfrtp_1 _24901_ (.CLK(clk_i),
    .D(_01749_),
    .RESET_B(net1559),
    .Q(\vmem[402] ));
 dfrtp_1 _24902_ (.CLK(clk_i),
    .D(_01750_),
    .RESET_B(net1555),
    .Q(\vmem[401] ));
 dfrtp_1 _24903_ (.CLK(clk_i),
    .D(_01751_),
    .RESET_B(net1517),
    .Q(\vmem[400] ));
 dfrtp_1 _24904_ (.CLK(clk_i),
    .D(_01752_),
    .RESET_B(net1534),
    .Q(\vmem[399] ));
 dfrtp_1 _24905_ (.CLK(clk_i),
    .D(_01753_),
    .RESET_B(net1546),
    .Q(\vmem[398] ));
 dfrtp_1 _24906_ (.CLK(clk_i),
    .D(_01754_),
    .RESET_B(net1541),
    .Q(\vmem[397] ));
 dfrtp_1 _24907_ (.CLK(clk_i),
    .D(_01755_),
    .RESET_B(net1566),
    .Q(\vmem[396] ));
 dfrtp_1 _24908_ (.CLK(clk_i),
    .D(_01756_),
    .RESET_B(net1543),
    .Q(\vmem[395] ));
 dfrtp_1 _24909_ (.CLK(clk_i),
    .D(_01757_),
    .RESET_B(net1519),
    .Q(\vmem[394] ));
 dfrtp_1 _24910_ (.CLK(clk_i),
    .D(_01758_),
    .RESET_B(net1549),
    .Q(\vmem[393] ));
 dfrtp_1 _24911_ (.CLK(clk_i),
    .D(_01759_),
    .RESET_B(net1519),
    .Q(\vmem[392] ));
 dfrtp_1 _24912_ (.CLK(clk_i),
    .D(_01760_),
    .RESET_B(net1524),
    .Q(\vmem[391] ));
 dfrtp_1 _24913_ (.CLK(clk_i),
    .D(_01761_),
    .RESET_B(net1572),
    .Q(\vmem[390] ));
 dfrtp_1 _24914_ (.CLK(clk_i),
    .D(_01762_),
    .RESET_B(net1518),
    .Q(\vmem[389] ));
 dfrtp_1 _24915_ (.CLK(clk_i),
    .D(_01763_),
    .RESET_B(net1562),
    .Q(\vmem[388] ));
 dfrtp_1 _24916_ (.CLK(clk_i),
    .D(_01764_),
    .RESET_B(net1510),
    .Q(\vmem[387] ));
 dfrtp_1 _24917_ (.CLK(clk_i),
    .D(_01765_),
    .RESET_B(net1559),
    .Q(\vmem[386] ));
 dfrtp_1 _24918_ (.CLK(clk_i),
    .D(_01766_),
    .RESET_B(net1567),
    .Q(\vmem[385] ));
 dfrtp_1 _24919_ (.CLK(clk_i),
    .D(_01767_),
    .RESET_B(net1527),
    .Q(\vmem[384] ));
 dfrtp_1 _24920_ (.CLK(clk_i),
    .D(_01768_),
    .RESET_B(net1532),
    .Q(\vmem[383] ));
 dfrtp_1 _24921_ (.CLK(clk_i),
    .D(_01769_),
    .RESET_B(net1543),
    .Q(\vmem[382] ));
 dfrtp_1 _24922_ (.CLK(clk_i),
    .D(_01770_),
    .RESET_B(net1540),
    .Q(\vmem[381] ));
 dfrtp_1 _24923_ (.CLK(clk_i),
    .D(_01771_),
    .RESET_B(net1576),
    .Q(\vmem[380] ));
 dfrtp_1 _24924_ (.CLK(clk_i),
    .D(_01772_),
    .RESET_B(net1536),
    .Q(\vmem[379] ));
 dfrtp_1 _24925_ (.CLK(clk_i),
    .D(_01773_),
    .RESET_B(net1522),
    .Q(\vmem[378] ));
 dfrtp_1 _24926_ (.CLK(clk_i),
    .D(_01774_),
    .RESET_B(net1549),
    .Q(\vmem[377] ));
 dfrtp_1 _24927_ (.CLK(clk_i),
    .D(_01775_),
    .RESET_B(net1521),
    .Q(\vmem[376] ));
 dfrtp_1 _24928_ (.CLK(clk_i),
    .D(_01776_),
    .RESET_B(net1529),
    .Q(\vmem[375] ));
 dfrtp_1 _24929_ (.CLK(clk_i),
    .D(_01777_),
    .RESET_B(net1576),
    .Q(\vmem[374] ));
 dfrtp_1 _24930_ (.CLK(clk_i),
    .D(_01778_),
    .RESET_B(net1508),
    .Q(\vmem[373] ));
 dfrtp_1 _24931_ (.CLK(clk_i),
    .D(_01779_),
    .RESET_B(net1562),
    .Q(\vmem[372] ));
 dfrtp_1 _24932_ (.CLK(clk_i),
    .D(_01780_),
    .RESET_B(net1506),
    .Q(\vmem[371] ));
 dfrtp_1 _24933_ (.CLK(clk_i),
    .D(_01781_),
    .RESET_B(net1551),
    .Q(\vmem[370] ));
 dfrtp_1 _24934_ (.CLK(clk_i),
    .D(_01782_),
    .RESET_B(net1551),
    .Q(\vmem[369] ));
 dfrtp_1 _24935_ (.CLK(clk_i),
    .D(_01783_),
    .RESET_B(net1526),
    .Q(\vmem[368] ));
 dfrtp_1 _24936_ (.CLK(clk_i),
    .D(_01784_),
    .RESET_B(net1532),
    .Q(\vmem[367] ));
 dfrtp_1 _24937_ (.CLK(clk_i),
    .D(_01785_),
    .RESET_B(net1546),
    .Q(\vmem[366] ));
 dfrtp_1 _24938_ (.CLK(clk_i),
    .D(_01786_),
    .RESET_B(net1540),
    .Q(\vmem[365] ));
 dfrtp_1 _24939_ (.CLK(clk_i),
    .D(_01787_),
    .RESET_B(net1576),
    .Q(\vmem[364] ));
 dfrtp_1 _24940_ (.CLK(clk_i),
    .D(_01788_),
    .RESET_B(net1538),
    .Q(\vmem[363] ));
 dfrtp_1 _24941_ (.CLK(clk_i),
    .D(_01789_),
    .RESET_B(net1522),
    .Q(\vmem[362] ));
 dfrtp_1 _24942_ (.CLK(clk_i),
    .D(_01790_),
    .RESET_B(net1549),
    .Q(\vmem[361] ));
 dfrtp_1 _24943_ (.CLK(clk_i),
    .D(_01791_),
    .RESET_B(net1521),
    .Q(\vmem[360] ));
 dfrtp_1 _24944_ (.CLK(clk_i),
    .D(_01792_),
    .RESET_B(net1529),
    .Q(\vmem[359] ));
 dfrtp_1 _24945_ (.CLK(clk_i),
    .D(_01793_),
    .RESET_B(net1577),
    .Q(\vmem[358] ));
 dfrtp_1 _24946_ (.CLK(clk_i),
    .D(_01794_),
    .RESET_B(net1512),
    .Q(\vmem[357] ));
 dfrtp_1 _24947_ (.CLK(clk_i),
    .D(_01795_),
    .RESET_B(net1570),
    .Q(\vmem[356] ));
 dfrtp_1 _24948_ (.CLK(clk_i),
    .D(_01796_),
    .RESET_B(net1507),
    .Q(\vmem[355] ));
 dfrtp_1 _24949_ (.CLK(clk_i),
    .D(_01797_),
    .RESET_B(net1552),
    .Q(\vmem[354] ));
 dfrtp_1 _24950_ (.CLK(clk_i),
    .D(_01798_),
    .RESET_B(net1554),
    .Q(\vmem[353] ));
 dfrtp_1 _24951_ (.CLK(clk_i),
    .D(_01799_),
    .RESET_B(net1526),
    .Q(\vmem[352] ));
 dfrtp_1 _24952_ (.CLK(clk_i),
    .D(_01800_),
    .RESET_B(net1535),
    .Q(\vmem[351] ));
 dfrtp_1 _24953_ (.CLK(clk_i),
    .D(_01801_),
    .RESET_B(net1544),
    .Q(\vmem[350] ));
 dfrtp_1 _24954_ (.CLK(clk_i),
    .D(_01802_),
    .RESET_B(net1540),
    .Q(\vmem[349] ));
 dfrtp_1 _24955_ (.CLK(clk_i),
    .D(_01803_),
    .RESET_B(net1576),
    .Q(\vmem[348] ));
 dfrtp_1 _24956_ (.CLK(clk_i),
    .D(_01804_),
    .RESET_B(net1538),
    .Q(\vmem[347] ));
 dfrtp_1 _24957_ (.CLK(clk_i),
    .D(_01805_),
    .RESET_B(net1523),
    .Q(\vmem[346] ));
 dfrtp_1 _24958_ (.CLK(clk_i),
    .D(_01806_),
    .RESET_B(net1549),
    .Q(\vmem[345] ));
 dfrtp_1 _24959_ (.CLK(clk_i),
    .D(_01807_),
    .RESET_B(net1520),
    .Q(\vmem[344] ));
 dfrtp_1 _24960_ (.CLK(clk_i),
    .D(_01808_),
    .RESET_B(net1524),
    .Q(\vmem[343] ));
 dfrtp_1 _24961_ (.CLK(clk_i),
    .D(_01809_),
    .RESET_B(net1571),
    .Q(\vmem[342] ));
 dfrtp_1 _24962_ (.CLK(clk_i),
    .D(_01810_),
    .RESET_B(net1512),
    .Q(\vmem[341] ));
 dfrtp_1 _24963_ (.CLK(clk_i),
    .D(_01811_),
    .RESET_B(net1562),
    .Q(\vmem[340] ));
 dfrtp_1 _24964_ (.CLK(clk_i),
    .D(_01812_),
    .RESET_B(net1510),
    .Q(\vmem[339] ));
 dfrtp_1 _24965_ (.CLK(clk_i),
    .D(_01813_),
    .RESET_B(net1558),
    .Q(\vmem[338] ));
 dfrtp_1 _24966_ (.CLK(clk_i),
    .D(_01814_),
    .RESET_B(net1565),
    .Q(\vmem[337] ));
 dfrtp_1 _24967_ (.CLK(clk_i),
    .D(_01815_),
    .RESET_B(net1526),
    .Q(\vmem[336] ));
 dfrtp_1 _24968_ (.CLK(clk_i),
    .D(_01816_),
    .RESET_B(net1532),
    .Q(\vmem[335] ));
 dfrtp_1 _24969_ (.CLK(clk_i),
    .D(_01817_),
    .RESET_B(net1544),
    .Q(\vmem[334] ));
 dfrtp_1 _24970_ (.CLK(clk_i),
    .D(_01818_),
    .RESET_B(net1540),
    .Q(\vmem[333] ));
 dfrtp_1 _24971_ (.CLK(clk_i),
    .D(_01819_),
    .RESET_B(net1576),
    .Q(\vmem[332] ));
 dfrtp_1 _24972_ (.CLK(clk_i),
    .D(_01820_),
    .RESET_B(net1536),
    .Q(\vmem[331] ));
 dfrtp_1 _24973_ (.CLK(clk_i),
    .D(_01821_),
    .RESET_B(net1523),
    .Q(\vmem[330] ));
 dfrtp_1 _24974_ (.CLK(clk_i),
    .D(_01822_),
    .RESET_B(net1528),
    .Q(\vmem[329] ));
 dfrtp_1 _24975_ (.CLK(clk_i),
    .D(_01823_),
    .RESET_B(net1519),
    .Q(\vmem[328] ));
 dfrtp_1 _24976_ (.CLK(clk_i),
    .D(_01824_),
    .RESET_B(net1524),
    .Q(\vmem[327] ));
 dfrtp_1 _24977_ (.CLK(clk_i),
    .D(_01825_),
    .RESET_B(net1577),
    .Q(\vmem[326] ));
 dfrtp_1 _24978_ (.CLK(clk_i),
    .D(_01826_),
    .RESET_B(net1513),
    .Q(\vmem[325] ));
 dfrtp_1 _24979_ (.CLK(clk_i),
    .D(_01827_),
    .RESET_B(net1563),
    .Q(\vmem[324] ));
 dfrtp_1 _24980_ (.CLK(clk_i),
    .D(_01828_),
    .RESET_B(net1510),
    .Q(\vmem[323] ));
 dfrtp_1 _24981_ (.CLK(clk_i),
    .D(_01829_),
    .RESET_B(net1558),
    .Q(\vmem[322] ));
 dfrtp_1 _24982_ (.CLK(clk_i),
    .D(_01830_),
    .RESET_B(net1565),
    .Q(\vmem[321] ));
 dfrtp_1 _24983_ (.CLK(clk_i),
    .D(_01831_),
    .RESET_B(net1526),
    .Q(\vmem[320] ));
 dfrtp_1 _24984_ (.CLK(clk_i),
    .D(_01832_),
    .RESET_B(net1535),
    .Q(\vmem[319] ));
 dfrtp_1 _24985_ (.CLK(clk_i),
    .D(_01833_),
    .RESET_B(net1544),
    .Q(\vmem[318] ));
 dfrtp_1 _24986_ (.CLK(clk_i),
    .D(_01834_),
    .RESET_B(net1540),
    .Q(\vmem[317] ));
 dfrtp_1 _24987_ (.CLK(clk_i),
    .D(_01835_),
    .RESET_B(net1568),
    .Q(\vmem[316] ));
 dfrtp_1 _24988_ (.CLK(clk_i),
    .D(_01836_),
    .RESET_B(net1536),
    .Q(\vmem[315] ));
 dfrtp_1 _24989_ (.CLK(clk_i),
    .D(_01837_),
    .RESET_B(net1525),
    .Q(\vmem[314] ));
 dfrtp_1 _24990_ (.CLK(clk_i),
    .D(_01838_),
    .RESET_B(net1549),
    .Q(\vmem[313] ));
 dfrtp_1 _24991_ (.CLK(clk_i),
    .D(_01839_),
    .RESET_B(net1521),
    .Q(\vmem[312] ));
 dfrtp_1 _24992_ (.CLK(clk_i),
    .D(_01840_),
    .RESET_B(net1528),
    .Q(\vmem[311] ));
 dfrtp_1 _24993_ (.CLK(clk_i),
    .D(_01841_),
    .RESET_B(net1571),
    .Q(\vmem[310] ));
 dfrtp_1 _24994_ (.CLK(clk_i),
    .D(_01842_),
    .RESET_B(net1515),
    .Q(\vmem[309] ));
 dfrtp_1 _24995_ (.CLK(clk_i),
    .D(_01843_),
    .RESET_B(net1563),
    .Q(\vmem[308] ));
 dfrtp_1 _24996_ (.CLK(clk_i),
    .D(_01844_),
    .RESET_B(net1507),
    .Q(\vmem[307] ));
 dfrtp_1 _24997_ (.CLK(clk_i),
    .D(_01845_),
    .RESET_B(net1549),
    .Q(\vmem[306] ));
 dfrtp_1 _24998_ (.CLK(clk_i),
    .D(_01846_),
    .RESET_B(net1554),
    .Q(\vmem[305] ));
 dfrtp_1 _24999_ (.CLK(clk_i),
    .D(_01847_),
    .RESET_B(net1526),
    .Q(\vmem[304] ));
 dfrtp_1 _25000_ (.CLK(clk_i),
    .D(_01848_),
    .RESET_B(net1532),
    .Q(\vmem[303] ));
 dfrtp_1 _25001_ (.CLK(clk_i),
    .D(_01849_),
    .RESET_B(net1546),
    .Q(\vmem[302] ));
 dfrtp_1 _25002_ (.CLK(clk_i),
    .D(_01850_),
    .RESET_B(net1542),
    .Q(\vmem[301] ));
 dfrtp_1 _25003_ (.CLK(clk_i),
    .D(_01851_),
    .RESET_B(net1568),
    .Q(\vmem[300] ));
 dfrtp_1 _25004_ (.CLK(clk_i),
    .D(_01852_),
    .RESET_B(net1536),
    .Q(\vmem[299] ));
 dfrtp_1 _25005_ (.CLK(clk_i),
    .D(_01853_),
    .RESET_B(net1523),
    .Q(\vmem[298] ));
 dfrtp_1 _25006_ (.CLK(clk_i),
    .D(_01854_),
    .RESET_B(net1550),
    .Q(\vmem[297] ));
 dfrtp_1 _25007_ (.CLK(clk_i),
    .D(_01855_),
    .RESET_B(net1521),
    .Q(\vmem[296] ));
 dfrtp_1 _25008_ (.CLK(clk_i),
    .D(_01856_),
    .RESET_B(net1550),
    .Q(\vmem[295] ));
 dfrtp_1 _25009_ (.CLK(clk_i),
    .D(_01857_),
    .RESET_B(net1571),
    .Q(\vmem[294] ));
 dfrtp_1 _25010_ (.CLK(clk_i),
    .D(_01858_),
    .RESET_B(net1515),
    .Q(\vmem[293] ));
 dfrtp_1 _25011_ (.CLK(clk_i),
    .D(_01859_),
    .RESET_B(net1570),
    .Q(\vmem[292] ));
 dfrtp_1 _25012_ (.CLK(clk_i),
    .D(_01860_),
    .RESET_B(net1507),
    .Q(\vmem[291] ));
 dfrtp_1 _25013_ (.CLK(clk_i),
    .D(_01861_),
    .RESET_B(net1550),
    .Q(\vmem[290] ));
 dfrtp_1 _25014_ (.CLK(clk_i),
    .D(_01862_),
    .RESET_B(net1554),
    .Q(\vmem[289] ));
 dfrtp_1 _25015_ (.CLK(clk_i),
    .D(_01863_),
    .RESET_B(net1527),
    .Q(\vmem[288] ));
 dfrtp_1 _25016_ (.CLK(clk_i),
    .D(_01864_),
    .RESET_B(net1535),
    .Q(\vmem[287] ));
 dfrtp_1 _25017_ (.CLK(clk_i),
    .D(_01865_),
    .RESET_B(net1544),
    .Q(\vmem[286] ));
 dfrtp_1 _25018_ (.CLK(clk_i),
    .D(_01866_),
    .RESET_B(net1543),
    .Q(\vmem[285] ));
 dfrtp_1 _25019_ (.CLK(clk_i),
    .D(_01867_),
    .RESET_B(net1571),
    .Q(\vmem[284] ));
 dfrtp_1 _25020_ (.CLK(clk_i),
    .D(_01868_),
    .RESET_B(net1536),
    .Q(\vmem[283] ));
 dfrtp_1 _25021_ (.CLK(clk_i),
    .D(_01869_),
    .RESET_B(net1525),
    .Q(\vmem[282] ));
 dfrtp_1 _25022_ (.CLK(clk_i),
    .D(_01870_),
    .RESET_B(net1528),
    .Q(\vmem[281] ));
 dfrtp_1 _25023_ (.CLK(clk_i),
    .D(_01871_),
    .RESET_B(net1519),
    .Q(\vmem[280] ));
 dfrtp_1 _25024_ (.CLK(clk_i),
    .D(_01872_),
    .RESET_B(net1529),
    .Q(\vmem[279] ));
 dfrtp_1 _25025_ (.CLK(clk_i),
    .D(_01873_),
    .RESET_B(net1571),
    .Q(\vmem[278] ));
 dfrtp_1 _25026_ (.CLK(clk_i),
    .D(_01874_),
    .RESET_B(net1515),
    .Q(\vmem[277] ));
 dfrtp_1 _25027_ (.CLK(clk_i),
    .D(_01875_),
    .RESET_B(net1563),
    .Q(\vmem[276] ));
 dfrtp_1 _25028_ (.CLK(clk_i),
    .D(_01876_),
    .RESET_B(net1510),
    .Q(\vmem[275] ));
 dfrtp_1 _25029_ (.CLK(clk_i),
    .D(_01877_),
    .RESET_B(net1556),
    .Q(\vmem[274] ));
 dfrtp_1 _25030_ (.CLK(clk_i),
    .D(_01878_),
    .RESET_B(net1555),
    .Q(\vmem[273] ));
 dfrtp_1 _25031_ (.CLK(clk_i),
    .D(_01879_),
    .RESET_B(net1515),
    .Q(\vmem[272] ));
 dfrtp_1 _25032_ (.CLK(clk_i),
    .D(_01880_),
    .RESET_B(net1532),
    .Q(\vmem[271] ));
 dfrtp_1 _25033_ (.CLK(clk_i),
    .D(_01881_),
    .RESET_B(net1544),
    .Q(\vmem[270] ));
 dfrtp_1 _25034_ (.CLK(clk_i),
    .D(_01882_),
    .RESET_B(net1542),
    .Q(\vmem[269] ));
 dfrtp_1 _25035_ (.CLK(clk_i),
    .D(_01883_),
    .RESET_B(net1571),
    .Q(\vmem[268] ));
 dfrtp_1 _25036_ (.CLK(clk_i),
    .D(_01884_),
    .RESET_B(net1536),
    .Q(\vmem[267] ));
 dfrtp_1 _25037_ (.CLK(clk_i),
    .D(_01885_),
    .RESET_B(net1523),
    .Q(\vmem[266] ));
 dfrtp_1 _25038_ (.CLK(clk_i),
    .D(_01886_),
    .RESET_B(net1550),
    .Q(\vmem[265] ));
 dfrtp_1 _25039_ (.CLK(clk_i),
    .D(_01887_),
    .RESET_B(net1548),
    .Q(\vmem[264] ));
 dfrtp_1 _25040_ (.CLK(clk_i),
    .D(_01888_),
    .RESET_B(net1529),
    .Q(\vmem[263] ));
 dfrtp_1 _25041_ (.CLK(clk_i),
    .D(_01889_),
    .RESET_B(net1571),
    .Q(\vmem[262] ));
 dfrtp_1 _25042_ (.CLK(clk_i),
    .D(_01890_),
    .RESET_B(net1515),
    .Q(\vmem[261] ));
 dfrtp_1 _25043_ (.CLK(clk_i),
    .D(_01891_),
    .RESET_B(net1563),
    .Q(\vmem[260] ));
 dfrtp_1 _25044_ (.CLK(clk_i),
    .D(_01892_),
    .RESET_B(net1510),
    .Q(\vmem[259] ));
 dfrtp_1 _25045_ (.CLK(clk_i),
    .D(_01893_),
    .RESET_B(net1558),
    .Q(\vmem[258] ));
 dfrtp_1 _25046_ (.CLK(clk_i),
    .D(_01894_),
    .RESET_B(net1565),
    .Q(\vmem[257] ));
 dfrtp_1 _25047_ (.CLK(clk_i),
    .D(_01895_),
    .RESET_B(net1516),
    .Q(\vmem[256] ));
 dfrtp_1 _25048_ (.CLK(clk_i),
    .D(_01896_),
    .RESET_B(net1533),
    .Q(\vmem[255] ));
 dfrtp_1 _25049_ (.CLK(clk_i),
    .D(_01897_),
    .RESET_B(net1546),
    .Q(\vmem[254] ));
 dfrtp_1 _25050_ (.CLK(clk_i),
    .D(_01898_),
    .RESET_B(net1560),
    .Q(\vmem[253] ));
 dfrtp_1 _25051_ (.CLK(clk_i),
    .D(_01899_),
    .RESET_B(net1567),
    .Q(\vmem[252] ));
 dfrtp_1 _25052_ (.CLK(clk_i),
    .D(_01900_),
    .RESET_B(net1535),
    .Q(\vmem[251] ));
 dfrtp_1 _25053_ (.CLK(clk_i),
    .D(_01901_),
    .RESET_B(net1520),
    .Q(\vmem[250] ));
 dfrtp_1 _25054_ (.CLK(clk_i),
    .D(_01902_),
    .RESET_B(net1528),
    .Q(\vmem[249] ));
 dfrtp_1 _25055_ (.CLK(clk_i),
    .D(_01903_),
    .RESET_B(net1511),
    .Q(\vmem[248] ));
 dfrtp_1 _25056_ (.CLK(clk_i),
    .D(_01904_),
    .RESET_B(net1528),
    .Q(\vmem[247] ));
 dfrtp_1 _25057_ (.CLK(clk_i),
    .D(_01905_),
    .RESET_B(net1569),
    .Q(\vmem[246] ));
 dfrtp_1 _25058_ (.CLK(clk_i),
    .D(_01906_),
    .RESET_B(net1509),
    .Q(\vmem[245] ));
 dfrtp_1 _25059_ (.CLK(clk_i),
    .D(_01907_),
    .RESET_B(net1561),
    .Q(\vmem[244] ));
 dfrtp_1 _25060_ (.CLK(clk_i),
    .D(_01908_),
    .RESET_B(net1505),
    .Q(\vmem[243] ));
 dfrtp_1 _25061_ (.CLK(clk_i),
    .D(_01909_),
    .RESET_B(net1558),
    .Q(\vmem[242] ));
 dfrtp_1 _25062_ (.CLK(clk_i),
    .D(_01910_),
    .RESET_B(net1554),
    .Q(\vmem[241] ));
 dfrtp_1 _25063_ (.CLK(clk_i),
    .D(_01911_),
    .RESET_B(net1515),
    .Q(\vmem[240] ));
 dfrtp_1 _25064_ (.CLK(clk_i),
    .D(_01912_),
    .RESET_B(net1531),
    .Q(\vmem[239] ));
 dfrtp_1 _25065_ (.CLK(clk_i),
    .D(_01913_),
    .RESET_B(net1545),
    .Q(\vmem[238] ));
 dfrtp_1 _25066_ (.CLK(clk_i),
    .D(_01914_),
    .RESET_B(net1556),
    .Q(\vmem[237] ));
 dfrtp_1 _25067_ (.CLK(clk_i),
    .D(_01915_),
    .RESET_B(net1567),
    .Q(\vmem[236] ));
 dfrtp_1 _25068_ (.CLK(clk_i),
    .D(_01916_),
    .RESET_B(net1537),
    .Q(\vmem[235] ));
 dfrtp_1 _25069_ (.CLK(clk_i),
    .D(_01917_),
    .RESET_B(net1520),
    .Q(\vmem[234] ));
 dfrtp_1 _25070_ (.CLK(clk_i),
    .D(_01918_),
    .RESET_B(net1549),
    .Q(\vmem[233] ));
 dfrtp_1 _25071_ (.CLK(clk_i),
    .D(_01919_),
    .RESET_B(net1511),
    .Q(\vmem[232] ));
 dfrtp_1 _25072_ (.CLK(clk_i),
    .D(_01920_),
    .RESET_B(net1528),
    .Q(\vmem[231] ));
 dfrtp_1 _25073_ (.CLK(clk_i),
    .D(_01921_),
    .RESET_B(net1569),
    .Q(\vmem[230] ));
 dfrtp_1 _25074_ (.CLK(clk_i),
    .D(_01922_),
    .RESET_B(net1509),
    .Q(\vmem[229] ));
 dfrtp_1 _25075_ (.CLK(clk_i),
    .D(_01923_),
    .RESET_B(net1563),
    .Q(\vmem[228] ));
 dfrtp_1 _25076_ (.CLK(clk_i),
    .D(_01924_),
    .RESET_B(net1506),
    .Q(\vmem[227] ));
 dfrtp_1 _25077_ (.CLK(clk_i),
    .D(_01925_),
    .RESET_B(net1558),
    .Q(\vmem[226] ));
 dfrtp_1 _25078_ (.CLK(clk_i),
    .D(_01926_),
    .RESET_B(net1555),
    .Q(\vmem[225] ));
 dfrtp_1 _25079_ (.CLK(clk_i),
    .D(_01927_),
    .RESET_B(net1515),
    .Q(\vmem[224] ));
 dfrtp_1 _25080_ (.CLK(clk_i),
    .D(_01928_),
    .RESET_B(net1533),
    .Q(\vmem[223] ));
 dfrtp_1 _25081_ (.CLK(clk_i),
    .D(_01929_),
    .RESET_B(net1543),
    .Q(\vmem[222] ));
 dfrtp_1 _25082_ (.CLK(clk_i),
    .D(_01930_),
    .RESET_B(net1545),
    .Q(\vmem[221] ));
 dfrtp_1 _25083_ (.CLK(clk_i),
    .D(_01931_),
    .RESET_B(net1565),
    .Q(\vmem[220] ));
 dfrtp_1 _25084_ (.CLK(clk_i),
    .D(_01932_),
    .RESET_B(net1537),
    .Q(\vmem[219] ));
 dfrtp_1 _25085_ (.CLK(clk_i),
    .D(_01933_),
    .RESET_B(net1522),
    .Q(\vmem[218] ));
 dfrtp_1 _25086_ (.CLK(clk_i),
    .D(_01934_),
    .RESET_B(net1527),
    .Q(\vmem[217] ));
 dfrtp_1 _25087_ (.CLK(clk_i),
    .D(_01935_),
    .RESET_B(net1510),
    .Q(\vmem[216] ));
 dfrtp_1 _25088_ (.CLK(clk_i),
    .D(_01936_),
    .RESET_B(net1528),
    .Q(\vmem[215] ));
 dfrtp_1 _25089_ (.CLK(clk_i),
    .D(_01937_),
    .RESET_B(net1569),
    .Q(\vmem[214] ));
 dfrtp_1 _25090_ (.CLK(clk_i),
    .D(_01938_),
    .RESET_B(net1510),
    .Q(\vmem[213] ));
 dfrtp_1 _25091_ (.CLK(clk_i),
    .D(_01939_),
    .RESET_B(net1561),
    .Q(\vmem[212] ));
 dfrtp_1 _25092_ (.CLK(clk_i),
    .D(_01940_),
    .RESET_B(net1505),
    .Q(\vmem[211] ));
 dfrtp_1 _25093_ (.CLK(clk_i),
    .D(_01941_),
    .RESET_B(net1558),
    .Q(\vmem[210] ));
 dfrtp_1 _25094_ (.CLK(clk_i),
    .D(_01942_),
    .RESET_B(net1554),
    .Q(\vmem[209] ));
 dfrtp_1 _25095_ (.CLK(clk_i),
    .D(_01943_),
    .RESET_B(net1515),
    .Q(\vmem[208] ));
 dfrtp_1 _25096_ (.CLK(clk_i),
    .D(_01944_),
    .RESET_B(net1533),
    .Q(\vmem[207] ));
 dfrtp_1 _25097_ (.CLK(clk_i),
    .D(_01945_),
    .RESET_B(net1545),
    .Q(\vmem[206] ));
 dfrtp_1 _25098_ (.CLK(clk_i),
    .D(_01946_),
    .RESET_B(net1541),
    .Q(\vmem[205] ));
 dfrtp_1 _25099_ (.CLK(clk_i),
    .D(_01947_),
    .RESET_B(net1566),
    .Q(\vmem[204] ));
 dfrtp_1 _25100_ (.CLK(clk_i),
    .D(_01948_),
    .RESET_B(net1537),
    .Q(\vmem[203] ));
 dfrtp_1 _25101_ (.CLK(clk_i),
    .D(_01949_),
    .RESET_B(net1520),
    .Q(\vmem[202] ));
 dfrtp_1 _25102_ (.CLK(clk_i),
    .D(_01950_),
    .RESET_B(net1527),
    .Q(\vmem[201] ));
 dfrtp_1 _25103_ (.CLK(clk_i),
    .D(_01951_),
    .RESET_B(net1510),
    .Q(\vmem[200] ));
 dfrtp_1 _25104_ (.CLK(clk_i),
    .D(_01952_),
    .RESET_B(net1528),
    .Q(\vmem[199] ));
 dfrtp_1 _25105_ (.CLK(clk_i),
    .D(_01953_),
    .RESET_B(net1569),
    .Q(\vmem[198] ));
 dfrtp_1 _25106_ (.CLK(clk_i),
    .D(_01954_),
    .RESET_B(net1513),
    .Q(\vmem[197] ));
 dfrtp_1 _25107_ (.CLK(clk_i),
    .D(_01955_),
    .RESET_B(net1560),
    .Q(\vmem[196] ));
 dfrtp_1 _25108_ (.CLK(clk_i),
    .D(_01956_),
    .RESET_B(net1505),
    .Q(\vmem[195] ));
 dfrtp_1 _25109_ (.CLK(clk_i),
    .D(_01957_),
    .RESET_B(net1565),
    .Q(\vmem[194] ));
 dfrtp_1 _25110_ (.CLK(clk_i),
    .D(_01958_),
    .RESET_B(net1555),
    .Q(\vmem[193] ));
 dfrtp_1 _25111_ (.CLK(clk_i),
    .D(_01959_),
    .RESET_B(net1515),
    .Q(\vmem[192] ));
 dfrtp_1 _25112_ (.CLK(clk_i),
    .D(_01960_),
    .RESET_B(net1533),
    .Q(\vmem[191] ));
 dfrtp_1 _25113_ (.CLK(clk_i),
    .D(_01961_),
    .RESET_B(net1545),
    .Q(\vmem[190] ));
 dfrtp_1 _25114_ (.CLK(clk_i),
    .D(_01962_),
    .RESET_B(net1541),
    .Q(\vmem[189] ));
 dfrtp_1 _25115_ (.CLK(clk_i),
    .D(_01963_),
    .RESET_B(net1565),
    .Q(\vmem[188] ));
 dfrtp_1 _25116_ (.CLK(clk_i),
    .D(_01964_),
    .RESET_B(net1537),
    .Q(\vmem[187] ));
 dfrtp_1 _25117_ (.CLK(clk_i),
    .D(_01965_),
    .RESET_B(net1520),
    .Q(\vmem[186] ));
 dfrtp_1 _25118_ (.CLK(clk_i),
    .D(_01966_),
    .RESET_B(net1553),
    .Q(\vmem[185] ));
 dfrtp_1 _25119_ (.CLK(clk_i),
    .D(_01967_),
    .RESET_B(net1511),
    .Q(\vmem[184] ));
 dfrtp_1 _25120_ (.CLK(clk_i),
    .D(_01968_),
    .RESET_B(net1528),
    .Q(\vmem[183] ));
 dfrtp_1 _25121_ (.CLK(clk_i),
    .D(_01969_),
    .RESET_B(net1569),
    .Q(\vmem[182] ));
 dfrtp_1 _25122_ (.CLK(clk_i),
    .D(_01970_),
    .RESET_B(net1512),
    .Q(\vmem[181] ));
 dfrtp_1 _25123_ (.CLK(clk_i),
    .D(_01971_),
    .RESET_B(net1561),
    .Q(\vmem[180] ));
 dfrtp_1 _25124_ (.CLK(clk_i),
    .D(_01972_),
    .RESET_B(net1506),
    .Q(\vmem[179] ));
 dfrtp_1 _25125_ (.CLK(clk_i),
    .D(_01973_),
    .RESET_B(net1556),
    .Q(\vmem[178] ));
 dfrtp_1 _25126_ (.CLK(clk_i),
    .D(_01974_),
    .RESET_B(net1578),
    .Q(\vmem[177] ));
 dfrtp_1 _25127_ (.CLK(clk_i),
    .D(_01975_),
    .RESET_B(net1517),
    .Q(\vmem[176] ));
 dfrtp_1 _25128_ (.CLK(clk_i),
    .D(_01976_),
    .RESET_B(net1531),
    .Q(\vmem[175] ));
 dfrtp_1 _25129_ (.CLK(clk_i),
    .D(_01977_),
    .RESET_B(net1560),
    .Q(\vmem[174] ));
 dfrtp_1 _25130_ (.CLK(clk_i),
    .D(_01978_),
    .RESET_B(net1557),
    .Q(\vmem[173] ));
 dfrtp_1 _25131_ (.CLK(clk_i),
    .D(_01979_),
    .RESET_B(net1565),
    .Q(\vmem[172] ));
 dfrtp_1 _25132_ (.CLK(clk_i),
    .D(_01980_),
    .RESET_B(net1537),
    .Q(\vmem[171] ));
 dfrtp_1 _25133_ (.CLK(clk_i),
    .D(_01981_),
    .RESET_B(net1520),
    .Q(\vmem[170] ));
 dfrtp_1 _25134_ (.CLK(clk_i),
    .D(_01982_),
    .RESET_B(net1553),
    .Q(\vmem[169] ));
 dfrtp_1 _25135_ (.CLK(clk_i),
    .D(_01983_),
    .RESET_B(net1511),
    .Q(\vmem[168] ));
 dfrtp_1 _25136_ (.CLK(clk_i),
    .D(_01984_),
    .RESET_B(net1530),
    .Q(\vmem[167] ));
 dfrtp_1 _25137_ (.CLK(clk_i),
    .D(_01985_),
    .RESET_B(net1571),
    .Q(\vmem[166] ));
 dfrtp_1 _25138_ (.CLK(clk_i),
    .D(_01986_),
    .RESET_B(net1512),
    .Q(\vmem[165] ));
 dfrtp_1 _25139_ (.CLK(clk_i),
    .D(_01987_),
    .RESET_B(net1563),
    .Q(\vmem[164] ));
 dfrtp_1 _25140_ (.CLK(clk_i),
    .D(_01988_),
    .RESET_B(net1506),
    .Q(\vmem[163] ));
 dfrtp_1 _25141_ (.CLK(clk_i),
    .D(_01989_),
    .RESET_B(net1550),
    .Q(\vmem[162] ));
 dfrtp_1 _25142_ (.CLK(clk_i),
    .D(_01990_),
    .RESET_B(net1578),
    .Q(\vmem[161] ));
 dfrtp_1 _25143_ (.CLK(clk_i),
    .D(_01991_),
    .RESET_B(net1517),
    .Q(\vmem[160] ));
 dfrtp_1 _25144_ (.CLK(clk_i),
    .D(_01992_),
    .RESET_B(net1533),
    .Q(\vmem[159] ));
 dfrtp_1 _25145_ (.CLK(clk_i),
    .D(_01993_),
    .RESET_B(net1545),
    .Q(\vmem[158] ));
 dfrtp_1 _25146_ (.CLK(clk_i),
    .D(_01994_),
    .RESET_B(net1541),
    .Q(\vmem[157] ));
 dfrtp_1 _25147_ (.CLK(clk_i),
    .D(_01995_),
    .RESET_B(net1566),
    .Q(\vmem[156] ));
 dfrtp_1 _25148_ (.CLK(clk_i),
    .D(_01996_),
    .RESET_B(net1537),
    .Q(\vmem[155] ));
 dfrtp_1 _25149_ (.CLK(clk_i),
    .D(_01997_),
    .RESET_B(net1520),
    .Q(\vmem[154] ));
 dfrtp_1 _25150_ (.CLK(clk_i),
    .D(_01998_),
    .RESET_B(net1553),
    .Q(\vmem[153] ));
 dfrtp_1 _25151_ (.CLK(clk_i),
    .D(_01999_),
    .RESET_B(net1510),
    .Q(\vmem[152] ));
 dfrtp_1 _25152_ (.CLK(clk_i),
    .D(_02000_),
    .RESET_B(net1530),
    .Q(\vmem[151] ));
 dfrtp_1 _25153_ (.CLK(clk_i),
    .D(_02001_),
    .RESET_B(net1569),
    .Q(\vmem[150] ));
 dfrtp_1 _25154_ (.CLK(clk_i),
    .D(_02002_),
    .RESET_B(net1510),
    .Q(\vmem[149] ));
 dfrtp_1 _25155_ (.CLK(clk_i),
    .D(_02003_),
    .RESET_B(net1561),
    .Q(\vmem[148] ));
 dfrtp_1 _25156_ (.CLK(clk_i),
    .D(_02004_),
    .RESET_B(net1506),
    .Q(\vmem[147] ));
 dfrtp_1 _25157_ (.CLK(clk_i),
    .D(_02005_),
    .RESET_B(net1556),
    .Q(\vmem[146] ));
 dfrtp_1 _25158_ (.CLK(clk_i),
    .D(_02006_),
    .RESET_B(net1555),
    .Q(\vmem[145] ));
 dfrtp_1 _25159_ (.CLK(clk_i),
    .D(_02007_),
    .RESET_B(net1517),
    .Q(\vmem[144] ));
 dfrtp_1 _25160_ (.CLK(clk_i),
    .D(_02008_),
    .RESET_B(net1533),
    .Q(\vmem[143] ));
 dfrtp_1 _25161_ (.CLK(clk_i),
    .D(_02009_),
    .RESET_B(net1545),
    .Q(\vmem[142] ));
 dfrtp_1 _25162_ (.CLK(clk_i),
    .D(_02010_),
    .RESET_B(net1542),
    .Q(\vmem[141] ));
 dfrtp_1 _25163_ (.CLK(clk_i),
    .D(_02011_),
    .RESET_B(net1566),
    .Q(\vmem[140] ));
 dfrtp_1 _25164_ (.CLK(clk_i),
    .D(_02012_),
    .RESET_B(net1537),
    .Q(\vmem[139] ));
 dfrtp_1 _25165_ (.CLK(clk_i),
    .D(_02013_),
    .RESET_B(net1520),
    .Q(\vmem[138] ));
 dfrtp_1 _25166_ (.CLK(clk_i),
    .D(_02014_),
    .RESET_B(net1527),
    .Q(\vmem[137] ));
 dfrtp_1 _25167_ (.CLK(clk_i),
    .D(_02015_),
    .RESET_B(net1511),
    .Q(\vmem[136] ));
 dfrtp_1 _25168_ (.CLK(clk_i),
    .D(_02016_),
    .RESET_B(net1528),
    .Q(\vmem[135] ));
 dfrtp_1 _25169_ (.CLK(clk_i),
    .D(_02017_),
    .RESET_B(net1571),
    .Q(\vmem[134] ));
 dfrtp_1 _25170_ (.CLK(clk_i),
    .D(_02018_),
    .RESET_B(net1512),
    .Q(\vmem[133] ));
 dfrtp_1 _25171_ (.CLK(clk_i),
    .D(_02019_),
    .RESET_B(net1561),
    .Q(\vmem[132] ));
 dfrtp_1 _25172_ (.CLK(clk_i),
    .D(_02020_),
    .RESET_B(net1506),
    .Q(\vmem[131] ));
 dfrtp_1 _25173_ (.CLK(clk_i),
    .D(_02021_),
    .RESET_B(net1556),
    .Q(\vmem[130] ));
 dfrtp_1 _25174_ (.CLK(clk_i),
    .D(_02022_),
    .RESET_B(net1555),
    .Q(\vmem[129] ));
 dfrtp_1 _25175_ (.CLK(clk_i),
    .D(_02023_),
    .RESET_B(net1517),
    .Q(\vmem[128] ));
 dfrtp_1 _25176_ (.CLK(clk_i),
    .D(_02024_),
    .RESET_B(net1531),
    .Q(\vmem[127] ));
 dfrtp_1 _25177_ (.CLK(clk_i),
    .D(_02025_),
    .RESET_B(net1543),
    .Q(\vmem[126] ));
 dfrtp_1 _25178_ (.CLK(clk_i),
    .D(_02026_),
    .RESET_B(net1540),
    .Q(\vmem[125] ));
 dfrtp_1 _25179_ (.CLK(clk_i),
    .D(_02027_),
    .RESET_B(net1576),
    .Q(\vmem[124] ));
 dfrtp_1 _25180_ (.CLK(clk_i),
    .D(_02028_),
    .RESET_B(net1535),
    .Q(\vmem[123] ));
 dfrtp_1 _25181_ (.CLK(clk_i),
    .D(_02029_),
    .RESET_B(net1522),
    .Q(\vmem[122] ));
 dfrtp_1 _25182_ (.CLK(clk_i),
    .D(_02030_),
    .RESET_B(net1551),
    .Q(\vmem[121] ));
 dfrtp_1 _25183_ (.CLK(clk_i),
    .D(_02031_),
    .RESET_B(net1519),
    .Q(\vmem[120] ));
 dfrtp_1 _25184_ (.CLK(clk_i),
    .D(_02032_),
    .RESET_B(net1529),
    .Q(\vmem[119] ));
 dfrtp_1 _25185_ (.CLK(clk_i),
    .D(_02033_),
    .RESET_B(net1577),
    .Q(\vmem[118] ));
 dfrtp_1 _25186_ (.CLK(clk_i),
    .D(_02034_),
    .RESET_B(net1508),
    .Q(\vmem[117] ));
 dfrtp_1 _25187_ (.CLK(clk_i),
    .D(_02035_),
    .RESET_B(net1562),
    .Q(\vmem[116] ));
 dfrtp_1 _25188_ (.CLK(clk_i),
    .D(_02036_),
    .RESET_B(net1505),
    .Q(\vmem[115] ));
 dfrtp_1 _25189_ (.CLK(clk_i),
    .D(_02037_),
    .RESET_B(net1557),
    .Q(\vmem[114] ));
 dfrtp_1 _25190_ (.CLK(clk_i),
    .D(_02038_),
    .RESET_B(net1554),
    .Q(\vmem[113] ));
 dfrtp_1 _25191_ (.CLK(clk_i),
    .D(_02039_),
    .RESET_B(net1517),
    .Q(\vmem[112] ));
 dfrtp_1 _25192_ (.CLK(clk_i),
    .D(_02040_),
    .RESET_B(net1531),
    .Q(\vmem[111] ));
 dfrtp_1 _25193_ (.CLK(clk_i),
    .D(_02041_),
    .RESET_B(net1545),
    .Q(\vmem[110] ));
 dfrtp_1 _25194_ (.CLK(clk_i),
    .D(_02042_),
    .RESET_B(net1542),
    .Q(\vmem[109] ));
 dfrtp_1 _25195_ (.CLK(clk_i),
    .D(_02043_),
    .RESET_B(net1576),
    .Q(\vmem[108] ));
 dfrtp_1 _25196_ (.CLK(clk_i),
    .D(_02044_),
    .RESET_B(net1535),
    .Q(\vmem[107] ));
 dfrtp_1 _25197_ (.CLK(clk_i),
    .D(_02045_),
    .RESET_B(net1522),
    .Q(\vmem[106] ));
 dfrtp_1 _25198_ (.CLK(clk_i),
    .D(_02046_),
    .RESET_B(net1553),
    .Q(\vmem[105] ));
 dfrtp_1 _25199_ (.CLK(clk_i),
    .D(_02047_),
    .RESET_B(net1519),
    .Q(\vmem[104] ));
 dfrtp_1 _25200_ (.CLK(clk_i),
    .D(_02048_),
    .RESET_B(net1529),
    .Q(\vmem[103] ));
 dfrtp_1 _25201_ (.CLK(clk_i),
    .D(_02049_),
    .RESET_B(net1577),
    .Q(\vmem[102] ));
 dfrtp_1 _25202_ (.CLK(clk_i),
    .D(_02050_),
    .RESET_B(net1508),
    .Q(\vmem[101] ));
 dfrtp_1 _25203_ (.CLK(clk_i),
    .D(_02051_),
    .RESET_B(net1569),
    .Q(\vmem[100] ));
 dfrtp_1 _25204_ (.CLK(clk_i),
    .D(_02052_),
    .RESET_B(net1506),
    .Q(\vmem[99] ));
 dfrtp_1 _25205_ (.CLK(clk_i),
    .D(_02053_),
    .RESET_B(net1556),
    .Q(\vmem[98] ));
 dfrtp_1 _25206_ (.CLK(clk_i),
    .D(_02054_),
    .RESET_B(net1554),
    .Q(\vmem[97] ));
 dfrtp_1 _25207_ (.CLK(clk_i),
    .D(_02055_),
    .RESET_B(net1517),
    .Q(\vmem[96] ));
 dfrtp_1 _25208_ (.CLK(clk_i),
    .D(_02056_),
    .RESET_B(net1531),
    .Q(\vmem[95] ));
 dfrtp_1 _25209_ (.CLK(clk_i),
    .D(_02057_),
    .RESET_B(net1543),
    .Q(\vmem[94] ));
 dfrtp_1 _25210_ (.CLK(clk_i),
    .D(_02058_),
    .RESET_B(net1540),
    .Q(\vmem[93] ));
 dfrtp_1 _25211_ (.CLK(clk_i),
    .D(_02059_),
    .RESET_B(net1576),
    .Q(\vmem[92] ));
 dfrtp_1 _25212_ (.CLK(clk_i),
    .D(_02060_),
    .RESET_B(net1535),
    .Q(\vmem[91] ));
 dfrtp_1 _25213_ (.CLK(clk_i),
    .D(_02061_),
    .RESET_B(net1523),
    .Q(\vmem[90] ));
 dfrtp_1 _25214_ (.CLK(clk_i),
    .D(_02062_),
    .RESET_B(net1553),
    .Q(\vmem[89] ));
 dfrtp_1 _25215_ (.CLK(clk_i),
    .D(_02063_),
    .RESET_B(net1519),
    .Q(\vmem[88] ));
 dfrtp_1 _25216_ (.CLK(clk_i),
    .D(_02064_),
    .RESET_B(net1525),
    .Q(\vmem[87] ));
 dfrtp_1 _25217_ (.CLK(clk_i),
    .D(_02065_),
    .RESET_B(net1572),
    .Q(\vmem[86] ));
 dfrtp_1 _25218_ (.CLK(clk_i),
    .D(_02066_),
    .RESET_B(net1509),
    .Q(\vmem[85] ));
 dfrtp_1 _25219_ (.CLK(clk_i),
    .D(_02067_),
    .RESET_B(net1563),
    .Q(\vmem[84] ));
 dfrtp_1 _25220_ (.CLK(clk_i),
    .D(_02068_),
    .RESET_B(net1505),
    .Q(\vmem[83] ));
 dfrtp_1 _25221_ (.CLK(clk_i),
    .D(_02069_),
    .RESET_B(net1557),
    .Q(\vmem[82] ));
 dfrtp_1 _25222_ (.CLK(clk_i),
    .D(_02070_),
    .RESET_B(net1552),
    .Q(\vmem[81] ));
 dfrtp_1 _25223_ (.CLK(clk_i),
    .D(_02071_),
    .RESET_B(net1516),
    .Q(\vmem[80] ));
 dfrtp_1 _25224_ (.CLK(clk_i),
    .D(_02072_),
    .RESET_B(net1531),
    .Q(\vmem[79] ));
 dfrtp_1 _25225_ (.CLK(clk_i),
    .D(_02073_),
    .RESET_B(net1543),
    .Q(\vmem[78] ));
 dfrtp_1 _25226_ (.CLK(clk_i),
    .D(_02074_),
    .RESET_B(net1533),
    .Q(\vmem[77] ));
 dfrtp_1 _25227_ (.CLK(clk_i),
    .D(_02075_),
    .RESET_B(net1576),
    .Q(\vmem[76] ));
 dfrtp_1 _25228_ (.CLK(clk_i),
    .D(_02076_),
    .RESET_B(net1535),
    .Q(\vmem[75] ));
 dfrtp_1 _25229_ (.CLK(clk_i),
    .D(_02077_),
    .RESET_B(net1522),
    .Q(\vmem[74] ));
 dfrtp_1 _25230_ (.CLK(clk_i),
    .D(_02078_),
    .RESET_B(net1553),
    .Q(\vmem[73] ));
 dfrtp_1 _25231_ (.CLK(clk_i),
    .D(_02079_),
    .RESET_B(net1511),
    .Q(\vmem[72] ));
 dfrtp_1 _25232_ (.CLK(clk_i),
    .D(_02080_),
    .RESET_B(net1524),
    .Q(\vmem[71] ));
 dfrtp_1 _25233_ (.CLK(clk_i),
    .D(_02081_),
    .RESET_B(net1577),
    .Q(\vmem[70] ));
 dfrtp_1 _25234_ (.CLK(clk_i),
    .D(_02082_),
    .RESET_B(net1509),
    .Q(\vmem[69] ));
 dfrtp_1 _25235_ (.CLK(clk_i),
    .D(_02083_),
    .RESET_B(net1562),
    .Q(\vmem[68] ));
 dfrtp_1 _25236_ (.CLK(clk_i),
    .D(_02084_),
    .RESET_B(net1505),
    .Q(\vmem[67] ));
 dfrtp_1 _25237_ (.CLK(clk_i),
    .D(_02085_),
    .RESET_B(net1557),
    .Q(\vmem[66] ));
 dfrtp_1 _25238_ (.CLK(clk_i),
    .D(_02086_),
    .RESET_B(net1554),
    .Q(\vmem[65] ));
 dfrtp_1 _25239_ (.CLK(clk_i),
    .D(_02087_),
    .RESET_B(net1516),
    .Q(\vmem[64] ));
 dfrtp_1 _25240_ (.CLK(clk_i),
    .D(_02088_),
    .RESET_B(net1531),
    .Q(\vmem[63] ));
 dfrtp_1 _25241_ (.CLK(clk_i),
    .D(_02089_),
    .RESET_B(net1560),
    .Q(\vmem[62] ));
 dfrtp_1 _25242_ (.CLK(clk_i),
    .D(_02090_),
    .RESET_B(net1542),
    .Q(\vmem[61] ));
 dfrtp_1 _25243_ (.CLK(clk_i),
    .D(_02091_),
    .RESET_B(net1567),
    .Q(\vmem[60] ));
 dfrtp_1 _25244_ (.CLK(clk_i),
    .D(_02092_),
    .RESET_B(net1536),
    .Q(\vmem[59] ));
 dfrtp_1 _25245_ (.CLK(clk_i),
    .D(_02093_),
    .RESET_B(net1524),
    .Q(\vmem[58] ));
 dfrtp_1 _25246_ (.CLK(clk_i),
    .D(_02094_),
    .RESET_B(net1549),
    .Q(\vmem[57] ));
 dfrtp_1 _25247_ (.CLK(clk_i),
    .D(_02095_),
    .RESET_B(net1519),
    .Q(\vmem[56] ));
 dfrtp_1 _25248_ (.CLK(clk_i),
    .D(_02096_),
    .RESET_B(net1529),
    .Q(\vmem[55] ));
 dfrtp_1 _25249_ (.CLK(clk_i),
    .D(_02097_),
    .RESET_B(net1572),
    .Q(\vmem[54] ));
 dfrtp_1 _25250_ (.CLK(clk_i),
    .D(_02098_),
    .RESET_B(net1508),
    .Q(\vmem[53] ));
 dfrtp_1 _25251_ (.CLK(clk_i),
    .D(_02099_),
    .RESET_B(net1562),
    .Q(\vmem[52] ));
 dfrtp_1 _25252_ (.CLK(clk_i),
    .D(_02100_),
    .RESET_B(net1508),
    .Q(\vmem[51] ));
 dfrtp_1 _25253_ (.CLK(clk_i),
    .D(_02101_),
    .RESET_B(net1558),
    .Q(\vmem[50] ));
 dfrtp_1 _25254_ (.CLK(clk_i),
    .D(_02102_),
    .RESET_B(net1551),
    .Q(\vmem[49] ));
 dfrtp_1 _25255_ (.CLK(clk_i),
    .D(_02103_),
    .RESET_B(net1516),
    .Q(\vmem[48] ));
 dfrtp_1 _25256_ (.CLK(clk_i),
    .D(_02104_),
    .RESET_B(net1531),
    .Q(\vmem[47] ));
 dfrtp_1 _25257_ (.CLK(clk_i),
    .D(_02105_),
    .RESET_B(net1560),
    .Q(\vmem[46] ));
 dfrtp_1 _25258_ (.CLK(clk_i),
    .D(_02106_),
    .RESET_B(net1542),
    .Q(\vmem[45] ));
 dfrtp_1 _25259_ (.CLK(clk_i),
    .D(_02107_),
    .RESET_B(net1567),
    .Q(\vmem[44] ));
 dfrtp_1 _25260_ (.CLK(clk_i),
    .D(_02108_),
    .RESET_B(net1536),
    .Q(\vmem[43] ));
 dfrtp_1 _25261_ (.CLK(clk_i),
    .D(_02109_),
    .RESET_B(net1522),
    .Q(\vmem[42] ));
 dfrtp_1 _25262_ (.CLK(clk_i),
    .D(_02110_),
    .RESET_B(net1549),
    .Q(\vmem[41] ));
 dfrtp_1 _25263_ (.CLK(clk_i),
    .D(_02111_),
    .RESET_B(net1519),
    .Q(\vmem[40] ));
 dfrtp_1 _25264_ (.CLK(clk_i),
    .D(_02112_),
    .RESET_B(net1529),
    .Q(\vmem[39] ));
 dfrtp_1 _25265_ (.CLK(clk_i),
    .D(_02113_),
    .RESET_B(net1572),
    .Q(\vmem[38] ));
 dfrtp_1 _25266_ (.CLK(clk_i),
    .D(_02114_),
    .RESET_B(net1508),
    .Q(\vmem[37] ));
 dfrtp_1 _25267_ (.CLK(clk_i),
    .D(_02115_),
    .RESET_B(net1569),
    .Q(\vmem[36] ));
 dfrtp_1 _25268_ (.CLK(clk_i),
    .D(_02116_),
    .RESET_B(net1508),
    .Q(\vmem[35] ));
 dfrtp_1 _25269_ (.CLK(clk_i),
    .D(_02117_),
    .RESET_B(net1557),
    .Q(\vmem[34] ));
 dfrtp_1 _25270_ (.CLK(clk_i),
    .D(_02118_),
    .RESET_B(net1554),
    .Q(\vmem[33] ));
 dfrtp_1 _25271_ (.CLK(clk_i),
    .D(_02119_),
    .RESET_B(net1515),
    .Q(\vmem[32] ));
 dfrtp_1 _25272_ (.CLK(clk_i),
    .D(_02120_),
    .RESET_B(net1531),
    .Q(\vmem[31] ));
 dfrtp_1 _25273_ (.CLK(clk_i),
    .D(_02121_),
    .RESET_B(net1543),
    .Q(\vmem[30] ));
 dfrtp_1 _25274_ (.CLK(clk_i),
    .D(_02122_),
    .RESET_B(net1541),
    .Q(\vmem[29] ));
 dfrtp_1 _25275_ (.CLK(clk_i),
    .D(_02123_),
    .RESET_B(net1567),
    .Q(\vmem[28] ));
 dfrtp_1 _25276_ (.CLK(clk_i),
    .D(_02124_),
    .RESET_B(net1535),
    .Q(\vmem[27] ));
 dfrtp_1 _25277_ (.CLK(clk_i),
    .D(_02125_),
    .RESET_B(net1522),
    .Q(\vmem[26] ));
 dfrtp_1 _25278_ (.CLK(clk_i),
    .D(_02126_),
    .RESET_B(net1553),
    .Q(\vmem[25] ));
 dfrtp_1 _25279_ (.CLK(clk_i),
    .D(_02127_),
    .RESET_B(net1520),
    .Q(\vmem[24] ));
 dfrtp_1 _25280_ (.CLK(clk_i),
    .D(_02128_),
    .RESET_B(net1525),
    .Q(\vmem[23] ));
 dfrtp_1 _25281_ (.CLK(clk_i),
    .D(_02129_),
    .RESET_B(net1572),
    .Q(\vmem[22] ));
 dfrtp_1 _25282_ (.CLK(clk_i),
    .D(_02130_),
    .RESET_B(net1509),
    .Q(\vmem[21] ));
 dfrtp_1 _25283_ (.CLK(clk_i),
    .D(_02131_),
    .RESET_B(net1562),
    .Q(\vmem[20] ));
 dfrtp_1 _25284_ (.CLK(clk_i),
    .D(_02132_),
    .RESET_B(net1505),
    .Q(\vmem[19] ));
 dfrtp_1 _25285_ (.CLK(clk_i),
    .D(_02133_),
    .RESET_B(net1557),
    .Q(\vmem[18] ));
 dfrtp_1 _25286_ (.CLK(clk_i),
    .D(_02134_),
    .RESET_B(net1552),
    .Q(\vmem[17] ));
 dfrtp_1 _25287_ (.CLK(clk_i),
    .D(_02135_),
    .RESET_B(net1516),
    .Q(\vmem[16] ));
 dfrtp_1 _25288_ (.CLK(clk_i),
    .D(_02136_),
    .RESET_B(net1532),
    .Q(\vmem[15] ));
 dfrtp_1 _25289_ (.CLK(clk_i),
    .D(_02137_),
    .RESET_B(net1543),
    .Q(\vmem[14] ));
 dfrtp_1 _25290_ (.CLK(clk_i),
    .D(_02138_),
    .RESET_B(net1540),
    .Q(\vmem[13] ));
 dfrtp_1 _25291_ (.CLK(clk_i),
    .D(_02139_),
    .RESET_B(net1568),
    .Q(\vmem[12] ));
 dfrtp_1 _25292_ (.CLK(clk_i),
    .D(_02140_),
    .RESET_B(net1535),
    .Q(\vmem[11] ));
 dfrtp_1 _25293_ (.CLK(clk_i),
    .D(_02141_),
    .RESET_B(net1522),
    .Q(\vmem[10] ));
 dfrtp_1 _25294_ (.CLK(clk_i),
    .D(_02142_),
    .RESET_B(net1553),
    .Q(\vmem[9] ));
 dfrtp_1 _25295_ (.CLK(clk_i),
    .D(_02143_),
    .RESET_B(net1519),
    .Q(\vmem[8] ));
 dfrtp_1 _25296_ (.CLK(clk_i),
    .D(_02144_),
    .RESET_B(net1524),
    .Q(\vmem[7] ));
 dfrtp_1 _25297_ (.CLK(clk_i),
    .D(_02145_),
    .RESET_B(net1572),
    .Q(\vmem[6] ));
 dfrtp_1 _25298_ (.CLK(clk_i),
    .D(_02146_),
    .RESET_B(net1509),
    .Q(\vmem[5] ));
 dfrtp_1 _25299_ (.CLK(clk_i),
    .D(_02147_),
    .RESET_B(net1562),
    .Q(\vmem[4] ));
 dfrtp_1 _25300_ (.CLK(clk_i),
    .D(_02148_),
    .RESET_B(net1575),
    .Q(\vmem[3] ));
 dfrtp_1 _25301_ (.CLK(clk_i),
    .D(_02149_),
    .RESET_B(net1559),
    .Q(\vmem[2] ));
 dfrtp_1 _25302_ (.CLK(clk_i),
    .D(_02150_),
    .RESET_B(net1554),
    .Q(\vmem[1] ));
 dfrtp_1 _25303_ (.CLK(clk_i),
    .D(_02151_),
    .RESET_B(net1516),
    .Q(\vmem[0] ));
 conb_1 _24009__1611 (.HI(net1611));
 conb_1 \digitop_pav2.rng_inst.rng_trngx_pav2.rngx_trngx_DONT_TOUCH.rngx_trngx_neg_data_DONT_TOUCH.stdinst_dfbbn_1_1612  (.HI(net1612));
 conb_1 \digitop_pav2.rng_inst.rng_trngx_pav2.rngx_trngx_DONT_TOUCH.rngx_trngx_neg_data_DONT_TOUCH.stdinst_dfbbn_1_1613  (.HI(net1613));
 conb_1 \digitop_pav2.sync_inst.inst_rstx.trigger_DONT_TOUCH1.stdinst_dfrtp_1_1614  (.HI(net1614));
 conb_1 \digitop_pav2.fm0miller_inst.fm0x_tx.muxdata_fmdata_0_1615  (.HI(net1615));
 conb_1 _24365__1583 (.LO(net1583));
 conb_1 _23621__1584 (.LO(net1584));
 conb_1 _23594__1585 (.LO(net1585));
 conb_1 \digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.stdinst_nor2_1_1586  (.LO(net1586));
 conb_1 \digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate1.stdinst_nor2_1_1587  (.LO(net1587));
 conb_1 \digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate2.stdinst_nor2_1_1588  (.LO(net1588));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gate.stdinst_nor2_1_1589  (.LO(net1589));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_gen_cg.stdinst_nor2_1_1590  (.LO(net1590));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_block_access.stdinst_nor2_1_1591  (.LO(net1591));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_block_ack.stdinst_nor2_1_1592  (.LO(net1592));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_block_invent.stdinst_nor2_1_1593  (.LO(net1593));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_block_sec.stdinst_nor2_1_1594  (.LO(net1594));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_boot.inst_gate.stdinst_nor2_1_1595  (.LO(net1595));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_cgate.stdinst_nor2_1_1596  (.LO(net1596));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_cipher.inst_gate.stdinst_nor2_1_1597  (.LO(net1597));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_gate.stdinst_nor2_1_1598  (.LO(net1598));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_fm0x.inst_gate.stdinst_nor2_1_1599  (.LO(net1599));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_gate.stdinst_or2_0_1600  (.LO(net1600));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.stdinst_nor2_1_1601  (.LO(net1601));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.stdinst_nor2_1_1602  (.LO(net1602));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.stdinst_nor2_1_1603  (.LO(net1603));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_gate.stdinst_nor2_1_1604  (.LO(net1604));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.stdinst_inv_1_1605  (.LO(net1605));
 conb_1 \digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.stdinst_nor2_1_1606  (.LO(net1606));
 conb_1 \digitop_pav2.sync_inst.inst_rstx.sync_rstx_gate.stdinst_nor2_1_1607  (.LO(net1607));
 conb_1 \digitop_pav2.fm0miller_inst.fm0x_tx.muxdata_fmdata_0_1608  (.LO(net1608));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_0.A ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_0.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_0.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_1.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_2.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_1.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_2.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_3.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_2.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_3.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_4.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_3.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_4.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_5.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_4.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_5.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_6.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_5.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_6.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_7.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_6.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_7.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_8.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_7.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_8.Y ));
 clkbuf_2 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_9.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_8.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b0_9.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_0.A ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_0.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_0.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_1.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_2.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_1.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_2.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_3.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_2.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_3.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_4.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_3.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_4.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_5.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_4.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_5.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_6.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_5.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_6.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_7.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_6.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_7.Y ));
 dlygate4sd3_1 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_8.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_7.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_8.Y ));
 buf_2 \digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_9.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_8.Y ),
    .X(\digitop_pav2.aes128_inst.stadly_aes128_counter_2b1_9.Y ));
 inv_1 \digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.stdinst_inv_1  (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.enable ),
    .Y(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.w_not ));
 nor2_1 \digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.stdinst_nor2_1  (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.w_not ),
    .B(net1586),
    .Y(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.w_nor ));
 or2_4 \digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.stdinst_or2_4  (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.w_nor ),
    .B(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.ck_in ),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.ck_out ));
 clkbuf_1 \digitop_pav2.cal_inst.dtest.calx_dtest_clk.sdcbuf_data_cgdis_stab_clk_is_data  (.A(_00133_),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.enable ));
 buf_2 \digitop_pav2.cal_inst.dtest.calx_dtest_clk.sdcbuf_dtest_auxclk  (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.aux_clk ),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.auxclk_after_buf ));
 buf_2 \digitop_pav2.cal_inst.dtest.calx_dtest_clk.sdcbuf_dtest_clk2  (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk2 ),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk2_after_buf ));
 buf_2 \digitop_pav2.cal_inst.dtest.calx_dtest_clk.sdcbuf_dtest_clk4  (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.clk4 ),
    .X(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.ck_in ));
 buf_2 \digitop_pav2.cal_inst.dtest.sdcbuf_stab_clk  (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.cal_stab_clk_cg.ck_out ),
    .X(\digitop_pav2.cal_inst.calx_clk_o ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[0].fm0miller_pav2_gand_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.gand ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[0].fm0miller_pav2_gand_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[0].fm0miller_pav2_gor_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[0].fm0miller_pav2_gor_dly.A ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[0].fm0miller_pav2_gor_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[1].fm0miller_pav2_gand_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[0].fm0miller_pav2_gand_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[1].fm0miller_pav2_gand_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[1].fm0miller_pav2_gor_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[0].fm0miller_pav2_gor_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[1].fm0miller_pav2_gor_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[2].fm0miller_pav2_gand_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[1].fm0miller_pav2_gand_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[2].fm0miller_pav2_gand_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[2].fm0miller_pav2_gor_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[1].fm0miller_pav2_gor_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[2].fm0miller_pav2_gor_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[3].fm0miller_pav2_gand_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[2].fm0miller_pav2_gand_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[3].fm0miller_pav2_gand_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[3].fm0miller_pav2_gor_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[2].fm0miller_pav2_gor_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[3].fm0miller_pav2_gor_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[4].fm0miller_pav2_gand_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[3].fm0miller_pav2_gand_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[4].fm0miller_pav2_gand_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[4].fm0miller_pav2_gor_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[3].fm0miller_pav2_gor_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[4].fm0miller_pav2_gor_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[5].fm0miller_pav2_gand_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[4].fm0miller_pav2_gand_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[5].fm0miller_pav2_gand_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[5].fm0miller_pav2_gor_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[4].fm0miller_pav2_gor_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[5].fm0miller_pav2_gor_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[6].fm0miller_pav2_gand_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[5].fm0miller_pav2_gand_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[6].fm0miller_pav2_gand_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[6].fm0miller_pav2_gor_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[5].fm0miller_pav2_gor_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[6].fm0miller_pav2_gor_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[7].fm0miller_pav2_gand_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[6].fm0miller_pav2_gand_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[7].fm0miller_pav2_gand_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[7].fm0miller_pav2_gor_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[6].fm0miller_pav2_gor_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[7].fm0miller_pav2_gor_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[8].fm0miller_pav2_gand_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[7].fm0miller_pav2_gand_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[8].fm0miller_pav2_gand_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[8].fm0miller_pav2_gor_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[7].fm0miller_pav2_gor_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[8].fm0miller_pav2_gor_dly.Y ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[9].fm0miller_pav2_gand_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[8].fm0miller_pav2_gand_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.gand_delay ));
 dlygate4sd3_1 \digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[9].fm0miller_pav2_gor_dly.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[8].fm0miller_pav2_gor_dly.Y ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.genblk1[9].fm0miller_pav2_gor_dly.Y ));
 conb_1 _24189__1610 (.HI(net1610));
 dlygate4sd3_1 hold1 (.A(net1631),
    .X(net1617));
 inv_1 \digitop_pav2.fm0miller_inst.fm0x_tx.inv_data_fm0x_clk_is_data  (.A(\digitop_pav2.fm0miller_inst.fm0x_tx.data_fm0x_clk_is_data_after_buf ),
    .Y(\digitop_pav2.fm0miller_inst.fm0x_tx.data_fm0x_clk_is_data_after_buf_b ));
 mux4_1 \digitop_pav2.fm0miller_inst.fm0x_tx.muxdata_fmdata_0  (.A0(net1608),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_tx.data_fm0x_clk_is_data_after_buf ),
    .A2(net1615),
    .A3(\digitop_pav2.fm0miller_inst.fm0x_tx.data_fm0x_clk_is_data_after_buf ),
    .S0(\digitop_pav2.fm0miller_inst.ctrl[0] ),
    .S1(\digitop_pav2.fm0miller_inst.ctrl[1] ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_tx.w_fmdata_mux_0 ));
 mux4_1 \digitop_pav2.fm0miller_inst.fm0x_tx.muxdata_fmdata_1  (.A0(\digitop_pav2.fm0miller_inst.fm0x_tx.data_fm0x_clk_is_data_after_buf_b ),
    .A1(net1616),
    .A2(\digitop_pav2.fm0miller_inst.fm0x_tx.data_fm0x_clk_is_data_after_buf_b ),
    .A3(net1609),
    .S0(\digitop_pav2.fm0miller_inst.ctrl[0] ),
    .S1(\digitop_pav2.fm0miller_inst.ctrl[1] ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_tx.w_fmdata_mux_1 ));
 mux2_1 \digitop_pav2.fm0miller_inst.fm0x_tx.muxdata_fmdata_2  (.A0(\digitop_pav2.fm0miller_inst.fm0x_tx.w_fmdata_mux_0 ),
    .A1(\digitop_pav2.fm0miller_inst.fm0x_tx.w_fmdata_mux_1 ),
    .S(\digitop_pav2.fm0miller_inst.ctrl[2] ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_mask.tx_raw_i ));
 buf_2 \digitop_pav2.fm0miller_inst.fm0x_tx.sdcbuf_data_fm0x_clk_is_data  (.A(\digitop_pav2.clkx_fm0x_clk ),
    .X(\digitop_pav2.fm0miller_inst.fm0x_tx.data_fm0x_clk_is_data_after_buf ));
 buf_2 \digitop_pav2.pie_inst.ctr.sdcbuf_pie_ctr_en  (.A(\digitop_pav2.pie_inst.ctr.en_ctr_i ),
    .X(\digitop_pav2.pie_inst.ctr.en_ctr_after_buf ));
 buf_2 \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.Y ));
 clkbuf_1 \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_1 \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[1].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_1 \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[2].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_1 \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[3].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_1 \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[4].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_1 \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[5].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_1 \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[6].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_1 \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[7].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_1 \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[8].piex_delay_buf1_DONT_TOUCH.Y ));
 buf_1 \digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.pie_inst.piex_ctr_clk_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_ctr_data_DONT_TOUCH.genblk1.genblk1.genblk1[9].piex_delay_buf1_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_en_ctr_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly1_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.en_ctr ),
    .X(\digitop_pav2.pie_inst.en_ctr_fix ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly1_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.clkx_irreg_clk ),
    .X(\digitop_pav2.pie_inst.fsm.clk_i ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly10_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly10_DONT_TOUCH.A ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly10_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly11_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly10_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly11_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly12_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly11_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly12_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly13_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly12_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly13_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly14_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly13_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly14_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly15_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly14_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly15_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly16_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly15_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly16_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly17_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly16_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly17_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly18_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly17_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly18_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly19_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly18_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly19_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly1_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.clkx_past_irreg_clk ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly1_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly20_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly19_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly20_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly21_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly20_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly21_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly22_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly21_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly22_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly23_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly22_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly23_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly24_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly23_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly24_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly25_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly24_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.fsm.past_clk_i ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly2_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly1_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly2_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly3_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly2_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly3_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly4_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly3_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly4_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly5_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly4_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly5_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly6_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly5_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly6_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly7_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly6_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly7_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly8_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly7_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly8_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly9_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly8_DONT_TOUCH.Y ),
    .X(\digitop_pav2.pie_inst.piex_past_irreg_clk_DONT_TOUCH.genblk1.genblk1.genblk1[0].piex_delay_dly10_DONT_TOUCH.A ));
 nor2_1 \digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate1.stdinst_nor2_1  (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.cg_en_out1 ),
    .B(net1587),
    .Y(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate1.w_nor ));
 or2_4 \digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate1.stdinst_or2_4  (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate1.w_nor ),
    .B(\digitop_pav2.clkx_cp_clk ),
    .X(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate1.ck_out ));
 nor2_1 \digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate2.stdinst_nor2_1  (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.cg_en_out2 ),
    .B(net1588),
    .Y(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate2.w_nor ));
 or2_4 \digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate2.stdinst_or2_4  (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate2.w_nor ),
    .B(\digitop_pav2.clkx_cp_clk ),
    .X(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_gate2.ck_out ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.blf_abort ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_0.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_0.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_1.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_2.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_1.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_2.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_3.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_2.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_3.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_4.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_3.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_4.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_5.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_4.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_5.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_6.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_5.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_6.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_7.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_6.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_7.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_8.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_7.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_8.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_9.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_8.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_blf_abort_9.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.dt_tx_st_o ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_0.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_0.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_1.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_2.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_1.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_2.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_3.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_2.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_3.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_4.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_3.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_4.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_5.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_4.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_5.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_6.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_5.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_6.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_7.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_6.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_7.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_8.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_7.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_8.Y ));
 buf_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_9.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_dt_tx_st_8.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.cmdfsm.fm0x_dt_tx_st_i ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.mod_en ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_0.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_0.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_1.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_2.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_1.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_2.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_3.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_2.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_3.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_4.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_3.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_4.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_5.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_4.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_5.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_6.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_5.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_6.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_7.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_6.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_7.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_8.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_7.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_8.Y ));
 clkbuf_2 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_9.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_fm0x_mod_en_8.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.cmdfsm.fm0x_mod_en_i ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmd_abort_b ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_0.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_0.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_1.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_2.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_1.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_2.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_3.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_2.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_3.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_4.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_3.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_4.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_5.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_4.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_5.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_6.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_5.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_6.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_7.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_6.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_7.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_8.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_7.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_8.Y ));
 clkbuf_1 \digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_9.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.stadly_proc_ctrl_pro_abort_b_8.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.cmdctr.pro_abort_b_i ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_0.stdinst_dlygate4sd3_1  (.A(net1302),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_0.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_0.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_1.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_2.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_1.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_2.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_3.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_2.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_3.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_4.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_3.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_4.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_5.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_4.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_5.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_6.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_5.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_6.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_7.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_6.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_7.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_8.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_7.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_8.Y ));
 dlymetal6s2s_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_9.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout2_DONT_TOUCH.stadly_proc_ctrl_int_8.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.ctr.piex_dt_rx_en_i ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.pass_t2_flag ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_0.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_0.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_1.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_2.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_1.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_2.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_3.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_2.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_3.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_4.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_3.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_4.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_5.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_4.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_5.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_6.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_5.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_6.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_7.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_6.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_7.Y ));
 dlygate4sd3_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_8.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_7.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_8.Y ));
 dlymetal6s2s_1 \digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_9.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.proc_ctrl_inst.timeout.proc_ctrl_timeout_DONT_TOUCH.stadly_proc_ctrl_int_8.Y ),
    .X(\digitop_pav2.proc_ctrl_inst.int_pass_t2_flag ));
 dfbbn_1 \digitop_pav2.rng_inst.rng_trngx_pav2.rngx_trngx_DONT_TOUCH.rngx_trngx_neg_data_DONT_TOUCH.stdinst_dfbbn_1  (.CLK_N(\digitop_pav2.clkx_rngx_clk ),
    .D(\digitop_pav2.clkx_rngx_fast_clk ),
    .RESET_B(net1612),
    .SET_B(net1613),
    .Q(\digitop_pav2.rng_inst.rng_trngx_pav2.neg_data ),
    .Q_N(\digitop_pav2.rng_inst.rng_trngx_pav2.rngx_trngx_DONT_TOUCH.neg_data_nc ));
 dfxtp_1 \digitop_pav2.rng_inst.rng_trngx_pav2.rngx_trngx_DONT_TOUCH.rngx_trngx_pos_data_DONT_TOUCH.stdinst_dfxtp_1  (.CLK(\digitop_pav2.clkx_rngx_clk ),
    .D(\digitop_pav2.clkx_rngx_fast_clk ),
    .Q(\digitop_pav2.rng_inst.rng_trngx_pav2.pos_data ));
 buf_2 \digitop_pav2.sdcbuf_fm0x_clk_for_proc_ctrl  (.A(\digitop_pav2.clkx_fm0x_clk ),
    .X(\digitop_pav2.fm0x_clk_for_proc_ctrl ));
 buf_2 \digitop_pav2.sdcbuf_func_clk  (.A(\digitop_pav2.func_clk_pre ),
    .X(\digitop_pav2.func_clk ));
 buf_2 \digitop_pav2.sdcbuf_s1_in  (.A(\digitop_pav2.s1_i ),
    .X(\digitop_pav2.invent_inst.s1_i ));
 clkbuf_4 \digitop_pav2.sdcbuf_s2_in  (.A(\digitop_pav2.s2_i ),
    .X(\digitop_pav2.invent_inst.invent_qqqr_pav2.s2_i ));
 clkbuf_4 \digitop_pav2.sdcbuf_s3_in  (.A(\digitop_pav2.s3_i ),
    .X(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ));
 clkbuf_4 \digitop_pav2.sdcbuf_sl_in  (.A(\digitop_pav2.sl_i ),
    .X(\digitop_pav2.invent_inst.invent_qqqr_pav2.sl_i ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_rd_en_0.stdinst_dlygate4sd3_1  (.A(net1705),
    .X(\digitop_pav2.stadly_memctrl_rd_en_0.Y ));
 clkbuf_2 \digitop_pav2.stadly_memctrl_rd_en_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_rd_en_0.Y ),
    .X(\digitop_pav2.memctrl_inst.nvm_rd_en_i ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt0_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt0_0.A ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt0_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt0_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt0_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt0_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt10_0.stdinst_dlygate4sd3_1  (.A(net1793),
    .X(\digitop_pav2.stadly_memctrl_wr_dt10_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt10_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt10_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt10_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt11_0.stdinst_dlygate4sd3_1  (.A(net1798),
    .X(\digitop_pav2.stadly_memctrl_wr_dt11_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt11_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt11_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt11_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt12_0.stdinst_dlygate4sd3_1  (.A(net1791),
    .X(\digitop_pav2.stadly_memctrl_wr_dt12_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt12_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt12_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt12_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt13_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt13_0.A ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt13_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt13_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt13_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt13_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt14_0.stdinst_dlygate4sd3_1  (.A(net1789),
    .X(\digitop_pav2.stadly_memctrl_wr_dt14_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt14_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt14_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt14_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt15_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt15_0.A ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt15_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt15_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt15_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt15_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt1_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt1_0.A ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt1_0.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt1_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt1_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt1_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt2_0.stdinst_dlygate4sd3_1  (.A(net1805),
    .X(\digitop_pav2.stadly_memctrl_wr_dt2_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt2_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt2_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt2_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt3_0.stdinst_dlygate4sd3_1  (.A(net1802),
    .X(\digitop_pav2.stadly_memctrl_wr_dt3_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt3_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt3_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt3_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt4_0.stdinst_dlygate4sd3_1  (.A(net1800),
    .X(\digitop_pav2.stadly_memctrl_wr_dt4_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt4_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt4_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt4_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt5_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt5_0.A ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt5_0.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt5_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt5_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt5_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt6_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt6_0.A ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt6_0.Y ));
 dlymetal6s2s_1 \digitop_pav2.stadly_memctrl_wr_dt6_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt6_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt6_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt7_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt7_0.A ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt7_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt7_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt7_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt7_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt8_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt8_0.A ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt8_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt8_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt8_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt8_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_dt9_0.stdinst_dlygate4sd3_1  (.A(net1796),
    .X(\digitop_pav2.stadly_memctrl_wr_dt9_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_dt9_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_dt9_0.Y ),
    .X(\digitop_pav2.stadly_memctrl_wr_dt9_1.Y ));
 dlygate4sd3_1 \digitop_pav2.stadly_memctrl_wr_en_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.glue_inst.mbus_wr_en_o ),
    .X(\digitop_pav2.stadly_memctrl_wr_en_0.Y ));
 buf_1 \digitop_pav2.stadly_memctrl_wr_en_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.stadly_memctrl_wr_en_0.Y ),
    .X(\digitop_pav2.memctrl_inst.nvm_wr_en_i ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 clkbuf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[5].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[5].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[5].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 buf_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[7].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[7].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[7].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[1].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[2].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[3].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[4].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[5].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[5].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[5].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_buf_2  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_blf_ctr_clk_DONT_TOUCH.genblk1.genblk1[6].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.sdcbuf_blf_ctr_rst_b  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_9.Y ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_0.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.rst_b_aux_before_buf ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_0.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_1.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_0.Y ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_1.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_2.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_1.Y ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_2.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_3.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_2.Y ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_3.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_4.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_3.Y ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_4.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_5.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_4.Y ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_5.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_6.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_5.Y ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_6.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_7.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_6.Y ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_7.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_8.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_7.Y ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_8.Y ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_9.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_8.Y ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_ctr.stadly_sync_blf_ctr_rst_b_9.Y ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.sdcbuf_mode_clk  (.A(net1250),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.mode_after_buf ));
 inv_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gate.stdinst_inv_1  (.A(\digitop_pav2.sync_inst.inst_clkx.en_blf_fc_b ),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gate.w_not ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gate.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gate.w_not ),
    .B(net1589),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gate.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gate.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gate.w_nor ),
    .B(\digitop_pav2.func_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_fc_clk_before_buf ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_gen_cg.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_gen_cg.enable ),
    .B(net1590),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_gen_cg.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_gen_cg.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_gen_cg.w_nor ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_fc_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_fc_clk_gated_before_buf ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.sdcbuf_blf_fc_clk_gated  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_fc_clk_gated_before_buf ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_gen.blf_fc_clk_gated ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.sdcbuf_blf_fc_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_fc_clk_before_buf ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_fc_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.sdcbuf_blf_pre_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_pre_clk_before_buf ),
    .X(\digitop_pav2.sync_inst.inst_clkx.blf_clk_pre ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.sdcbuf_blf_raw_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk_before_buf ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_blf.sdcbuf_blf_raw_mask  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_mask_before_buf ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_blf.blf_raw_mask ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_block_access.stdinst_nor2_1  (.A(net1194),
    .B(net1591),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_block_access.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_block_access.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_block_access.w_nor ),
    .B(\digitop_pav2.clkx_cp_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.access_clk_before_buf ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_block_ack.stdinst_nor2_1  (.A(net1266),
    .B(net1592),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_block_ack.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_block_ack.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_block_ack.w_nor ),
    .B(\digitop_pav2.clkx_cp_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.ack_clk_before_buf ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_block_invent.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.g_invent ),
    .B(net1593),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_block_invent.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_block_invent.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_block_invent.w_nor ),
    .B(\digitop_pav2.clkx_cp_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_block_invent.ck_out ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_block_sec.stdinst_nor2_1  (.A(net1004),
    .B(net1594),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_block_sec.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_block_sec.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_block_sec.w_nor ),
    .B(\digitop_pav2.clkx_cp_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_block_sec.ck_out ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_boot.inst_boot_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.boot_inst.r_boot_ff ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_boot.boot_dis_fix ));
 inv_1 \digitop_pav2.sync_inst.inst_clkx.inst_boot.inst_gate.stdinst_inv_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_boot.boot_dis_fix ),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_boot.inst_gate.w_not ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_boot.inst_gate.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_boot.inst_gate.w_not ),
    .B(net1595),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_boot.inst_gate.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_boot.inst_gate.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_boot.inst_gate.w_nor ),
    .B(\digitop_pav2.sync_inst.inst_clkx.dft_div4_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.boot_clk_before_buf ));
 inv_1 \digitop_pav2.sync_inst.inst_clkx.inst_cgate.stdinst_inv_1  (.A(\digitop_pav2.aes128_inst.aes128_regs.aes_exe_o ),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_cgate.w_not ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_cgate.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cgate.w_not ),
    .B(net1596),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_cgate.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_cgate.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cgate.w_nor ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_cgate.ck_in ),
    .X(\digitop_pav2.sync_inst.inst_clkx.blf_clk_before_buf ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_cipher.inst_gate.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cipher.cipher_en ),
    .B(net1597),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_cipher.inst_gate.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_cipher.inst_gate.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cipher.inst_gate.w_nor ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_cgate.ck_in ),
    .X(\digitop_pav2.sync_inst.inst_clkx.cipher_clk_before_buf ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_cp.auxbuf_cp  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_before_buf ),
    .X(\digitop_pav2.clkx_cp_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_cp.auxbuf_cp_div  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.div_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_div_after_buf ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_cp.auxbuf_cp_div_sel_0  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.cp_div_sel[0] ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.cp_div_sel_0_after_buf ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_cp.auxbuf_cp_div_sel_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.cp_div_sel[1] ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.cp_div_sel_1_after_buf ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_cp.auxbuf_cp_irreg  (.A(\digitop_pav2.clkx_irreg_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_irreg_after_buf ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_cp.auxbuf_cp_mode  (.A(net1250),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_mode_after_buf ));
 mux2_1 \digitop_pav2.sync_inst.inst_clkx.inst_cp.sdcbuf_cp_clk  (.A0(\digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_irreg_after_buf ),
    .A1(\digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_div_after_buf ),
    .S(\digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_mode_after_buf ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.aux_cp_before_buf ));
 mux4_1 \digitop_pav2.sync_inst.inst_clkx.inst_cp.sdcbuf_cp_div_clk  (.A0(\digitop_pav2.sync_inst.inst_clkx.blf_clk ),
    .A1(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m2_clk_after_buf ),
    .A2(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m4_clk_after_buf ),
    .A3(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m8_clk_after_buf ),
    .S0(\digitop_pav2.sync_inst.inst_clkx.inst_cp.cp_div_sel_0_after_buf ),
    .S1(\digitop_pav2.sync_inst.inst_clkx.inst_cp.cp_div_sel_1_after_buf ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.div_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_cp.sdcbuf_m2_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m2_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m2_clk_after_buf ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_cp.sdcbuf_m4_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m4_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m4_clk_after_buf ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_cp.sdcbuf_m8_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m8_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cp.m8_clk_after_buf ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.sdcbuf_div2_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.div2 ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.div2_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.sdcbuf_div4_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div.div4 ),
    .X(\digitop_pav2.sync_inst.inst_clkx.dft_div4_clk ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div4_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div4_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div4_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 inv_1 \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_gate.stdinst_inv_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_div4_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_gate.w_not ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_gate.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_gate.w_not ),
    .B(net1598),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_gate.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_gate.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_div4.inst_gate.w_nor ),
    .B(\digitop_pav2.func_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_div4.div_gated_clk_before_buf ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_div4.sdcbuf_div_gated_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_div4.div_gated_clk_before_buf ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_div4.div_gated_clk ));
 inv_1 \digitop_pav2.sync_inst.inst_clkx.inst_fm0x.inst_gate.stdinst_inv_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_fm0x.en_fm0x_clk_b ),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_fm0x.inst_gate.w_not ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_fm0x.inst_gate.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_fm0x.inst_gate.w_not ),
    .B(net1599),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_fm0x.inst_gate.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_fm0x.inst_gate.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_fm0x.inst_gate.w_nor ),
    .B(\digitop_pav2.sync_inst.inst_clkx.blf_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.fm0x_clk_before_buf ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_irreg.sdcbuf_pie_ff2_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_ff2 ),
    .X(\digitop_pav2.clkx_past_irreg_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_irreg.sdcbuf_pie_ff3_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_ff3 ),
    .X(\digitop_pav2.clkx_irreg_clk ));
 and2_4 \digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_gate.stdinst_and2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_gate.w_or ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_en.merge_clk_i ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_gate.ck_out ));
 or2_0 \digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_gate.stdinst_or2_0  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_mem.en_mem_clk ),
    .B(net1600),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_gate.w_or ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_mem.sdcbuf_mem_merge_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_merge.merge_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_en.merge_clk_i ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_mem.sdcbuf_mem_top_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_mem.inst_gate.ck_out ),
    .X(\digitop_pav2.clkx_mem_top_clk ));
 inv_1 \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.stdinst_inv_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.enable ),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.w_not ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.w_not ),
    .B(net1601),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.w_nor ),
    .B(\digitop_pav2.func_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_piex.clkx_piex_clk_o ));
 dlygate4sd3_1 \digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_piex_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_en.piex_clk_dis ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_piex.inst_gate.enable ));
 inv_1 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.stdinst_inv_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.en_pup_clk_b ),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.w_not ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.w_not ),
    .B(net1602),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.w_nor ),
    .B(\digitop_pav2.func_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.ck_out ));
 inv_1 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.stdinst_inv_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.en_pup_clk_b ),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.w_not ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.w_not ),
    .B(net1603),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.w_nor ),
    .B(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.scwend_clk_i ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.ck_out ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_rngx_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.slow_clk_en ),
    .X(\digitop_pav2.func_rnclk_en ));
 inv_1 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_gate.stdinst_inv_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.en_scwend_clk_b ),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_gate.w_not ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_gate.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_gate.w_not ),
    .B(net1604),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_gate.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_gate.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_gate.w_nor ),
    .B(rnclk_i),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.sdcbuf_boot_dis_clk  (.A(\digitop_pav2.boot_inst.r_boot_ff ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.boot_dis_clk_after_buf ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.sdcbuf_rngx_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_sel.rngx_clk ),
    .X(\digitop_pav2.clkx_rngx_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.sdcbuf_rngx_fast_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate0.ck_out ),
    .X(\digitop_pav2.clkx_rngx_fast_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.sdcbuf_rngx_pup_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_gate1.ck_out ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.rngx_pup_clk_i ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.sdcbuf_scwend_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_scwend.scwend_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.scwend_clk_i ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_rngx.sdcbuf_trigger_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_trigger.trigger_clk ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.trigger_clk_i ));
 inv_1 \digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.stdinst_inv_1  (.A(net1605),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.w_not ));
 nor2_1 \digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.w_not ),
    .B(net1606),
    .Y(\digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.w_nor ),
    .B(\digitop_pav2.sync_inst.inst_clkx.blf_clk_pre ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.ck_out ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.inst_wgate.sdcbuf_wgate_blf_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_wgate.inst_gate.ck_out ),
    .X(\digitop_pav2.sync_inst.inst_clkx.inst_cgate.ck_in ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.sdcbuf_access_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.access_clk_before_buf ),
    .X(\digitop_pav2.access_inst.access_check0.clk_i ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.sdcbuf_ack_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.ack_clk_before_buf ),
    .X(\digitop_pav2.ack_inst.clk_i ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.sdcbuf_blf_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.blf_clk_before_buf ),
    .X(\digitop_pav2.sync_inst.inst_clkx.blf_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.sdcbuf_boot_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.boot_clk_before_buf ),
    .X(\digitop_pav2.boot_inst.boot_ctrl0.clk_i ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.sdcbuf_cipher_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.cipher_clk_before_buf ),
    .X(\digitop_pav2.aes128_inst.aes128_counter.clk_i ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.sdcbuf_fm0x_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.fm0x_clk_before_buf ),
    .X(\digitop_pav2.clkx_fm0x_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.sdcbuf_invent_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_block_invent.ck_out ),
    .X(\digitop_pav2.clkx_invent_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.sdcbuf_piex_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_piex.clkx_piex_clk_o ),
    .X(\digitop_pav2.clkx_piex_clk ));
 buf_2 \digitop_pav2.sync_inst.inst_clkx.sdcbuf_sec_clk  (.A(\digitop_pav2.sync_inst.inst_clkx.inst_block_sec.ck_out ),
    .X(\digitop_pav2.clkx_sec_clk ));
 dlymetal6s2s_1 \digitop_pav2.sync_inst.inst_rstx.sync_rstx_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.stdinst_dlygate4sd3_1  (.A(net1825),
    .X(\digitop_pav2.sync_inst.inst_rstx.sync_rstx_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.Y ));
 inv_1 \digitop_pav2.sync_inst.inst_rstx.sync_rstx_gate.stdinst_inv_1  (.A(net1446),
    .Y(\digitop_pav2.sync_inst.inst_rstx.sync_rstx_gate.w_not ));
 nor2_1 \digitop_pav2.sync_inst.inst_rstx.sync_rstx_gate.stdinst_nor2_1  (.A(\digitop_pav2.sync_inst.inst_rstx.sync_rstx_gate.w_not ),
    .B(net1607),
    .Y(\digitop_pav2.sync_inst.inst_rstx.sync_rstx_gate.w_nor ));
 or2_4 \digitop_pav2.sync_inst.inst_rstx.sync_rstx_gate.stdinst_or2_4  (.A(\digitop_pav2.sync_inst.inst_rstx.sync_rstx_gate.w_nor ),
    .B(\digitop_pav2.func_clk ),
    .X(\digitop_pav2.sync_inst.inst_rstx.osc_clk_gated ));
 dfrtp_1 \digitop_pav2.sync_inst.inst_rstx.trigger_DONT_TOUCH1.stdinst_dfrtp_1  (.CLK(\digitop_pav2.sync_inst.inst_rstx.osc_clk_gated ),
    .D(net1614),
    .RESET_B(net1581),
    .Q(\digitop_pav2.sync_inst.inst_rstx.trigger_DONT_TOUCH1.Q ));
 dfrtp_1 \digitop_pav2.sync_inst.inst_rstx.trigger_DONT_TOUCH2.stdinst_dfrtp_1  (.CLK(\digitop_pav2.sync_inst.inst_rstx.osc_clk_gated ),
    .D(net1839),
    .RESET_B(net1581),
    .Q(\digitop_pav2.sync_inst.inst_rstx.sync_rstx_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ));
 buf_2 \digitop_pav2.testctrl_pav2.inst_enter.sdcbuf_tmrboot_clk  (.A(\digitop_pav2.boot_inst.r_boot_ff ),
    .X(\digitop_pav2.testctrl_pav2.inst_enter.tmrboot_clk ));
 and2_1 \digitop_pav2.testctrl_pav2.inst_tmamux.inst_and_sel_ibias  (.A(\digitop_pav2.testctrl_pav2.inst_tmamux.window_ibias ),
    .B(\digitop_pav2.testctrl_pav2.inst_tmamux.data_tclk_is_data ),
    .X(net71));
 and2_1 \digitop_pav2.testctrl_pav2.inst_tmamux.inst_and_sel_vcc  (.A(\digitop_pav2.testctrl_pav2.inst_tmamux.window_vcc ),
    .B(\digitop_pav2.testctrl_pav2.inst_tmamux.data_tclk_is_data ),
    .X(net72));
 and2_1 \digitop_pav2.testctrl_pav2.inst_tmamux.inst_and_sel_vdd  (.A(\digitop_pav2.testctrl_pav2.inst_tmamux.window_vdd ),
    .B(\digitop_pav2.testctrl_pav2.inst_tmamux.data_tclk_is_data ),
    .X(net73));
 and2_1 \digitop_pav2.testctrl_pav2.inst_tmamux.inst_and_sel_vref  (.A(\digitop_pav2.testctrl_pav2.inst_tmamux.window_vref ),
    .B(\digitop_pav2.testctrl_pav2.inst_tmamux.data_tclk_is_data ),
    .X(net74));
 buf_2 \digitop_pav2.testctrl_pav2.inst_tmamux.sdcbuf_data_tclk_is_data  (.A(tclk_i),
    .X(\digitop_pav2.testctrl_pav2.inst_tmamux.data_tclk_is_data ));
 clkbuf_1 \gen_obs_vmem[0].sdcbuf_gen_vmem  (.A(\vmem[0] ),
    .X(\vmem_after_buf[0] ));
 clkbuf_1 \gen_obs_vmem[100].sdcbuf_gen_vmem  (.A(\vmem[100] ),
    .X(\vmem_after_buf[100] ));
 clkbuf_1 \gen_obs_vmem[101].sdcbuf_gen_vmem  (.A(\vmem[101] ),
    .X(\vmem_after_buf[101] ));
 clkbuf_1 \gen_obs_vmem[102].sdcbuf_gen_vmem  (.A(\vmem[102] ),
    .X(\vmem_after_buf[102] ));
 clkbuf_1 \gen_obs_vmem[103].sdcbuf_gen_vmem  (.A(\vmem[103] ),
    .X(\vmem_after_buf[103] ));
 clkbuf_1 \gen_obs_vmem[104].sdcbuf_gen_vmem  (.A(\vmem[104] ),
    .X(\vmem_after_buf[104] ));
 clkbuf_1 \gen_obs_vmem[105].sdcbuf_gen_vmem  (.A(\vmem[105] ),
    .X(\vmem_after_buf[105] ));
 clkbuf_1 \gen_obs_vmem[106].sdcbuf_gen_vmem  (.A(\vmem[106] ),
    .X(\vmem_after_buf[106] ));
 clkbuf_1 \gen_obs_vmem[107].sdcbuf_gen_vmem  (.A(\vmem[107] ),
    .X(\vmem_after_buf[107] ));
 clkbuf_1 \gen_obs_vmem[108].sdcbuf_gen_vmem  (.A(\vmem[108] ),
    .X(\vmem_after_buf[108] ));
 clkbuf_1 \gen_obs_vmem[109].sdcbuf_gen_vmem  (.A(\vmem[109] ),
    .X(\vmem_after_buf[109] ));
 clkbuf_1 \gen_obs_vmem[10].sdcbuf_gen_vmem  (.A(\vmem[10] ),
    .X(\vmem_after_buf[10] ));
 clkbuf_1 \gen_obs_vmem[110].sdcbuf_gen_vmem  (.A(\vmem[110] ),
    .X(\vmem_after_buf[110] ));
 clkbuf_1 \gen_obs_vmem[111].sdcbuf_gen_vmem  (.A(\vmem[111] ),
    .X(\vmem_after_buf[111] ));
 clkbuf_1 \gen_obs_vmem[112].sdcbuf_gen_vmem  (.A(\vmem[112] ),
    .X(\vmem_after_buf[112] ));
 clkbuf_1 \gen_obs_vmem[113].sdcbuf_gen_vmem  (.A(\vmem[113] ),
    .X(\vmem_after_buf[113] ));
 clkbuf_1 \gen_obs_vmem[114].sdcbuf_gen_vmem  (.A(\vmem[114] ),
    .X(\vmem_after_buf[114] ));
 clkbuf_1 \gen_obs_vmem[115].sdcbuf_gen_vmem  (.A(\vmem[115] ),
    .X(\vmem_after_buf[115] ));
 clkbuf_1 \gen_obs_vmem[116].sdcbuf_gen_vmem  (.A(\vmem[116] ),
    .X(\vmem_after_buf[116] ));
 clkbuf_1 \gen_obs_vmem[117].sdcbuf_gen_vmem  (.A(\vmem[117] ),
    .X(\vmem_after_buf[117] ));
 clkbuf_1 \gen_obs_vmem[118].sdcbuf_gen_vmem  (.A(\vmem[118] ),
    .X(\vmem_after_buf[118] ));
 clkbuf_1 \gen_obs_vmem[119].sdcbuf_gen_vmem  (.A(\vmem[119] ),
    .X(\vmem_after_buf[119] ));
 clkbuf_1 \gen_obs_vmem[11].sdcbuf_gen_vmem  (.A(\vmem[11] ),
    .X(\vmem_after_buf[11] ));
 clkbuf_1 \gen_obs_vmem[120].sdcbuf_gen_vmem  (.A(\vmem[120] ),
    .X(\vmem_after_buf[120] ));
 clkbuf_1 \gen_obs_vmem[121].sdcbuf_gen_vmem  (.A(\vmem[121] ),
    .X(\vmem_after_buf[121] ));
 clkbuf_1 \gen_obs_vmem[122].sdcbuf_gen_vmem  (.A(\vmem[122] ),
    .X(\vmem_after_buf[122] ));
 clkbuf_1 \gen_obs_vmem[123].sdcbuf_gen_vmem  (.A(\vmem[123] ),
    .X(\vmem_after_buf[123] ));
 clkbuf_1 \gen_obs_vmem[124].sdcbuf_gen_vmem  (.A(\vmem[124] ),
    .X(\vmem_after_buf[124] ));
 clkbuf_1 \gen_obs_vmem[125].sdcbuf_gen_vmem  (.A(\vmem[125] ),
    .X(\vmem_after_buf[125] ));
 clkbuf_1 \gen_obs_vmem[126].sdcbuf_gen_vmem  (.A(\vmem[126] ),
    .X(\vmem_after_buf[126] ));
 clkbuf_1 \gen_obs_vmem[127].sdcbuf_gen_vmem  (.A(\vmem[127] ),
    .X(\vmem_after_buf[127] ));
 clkbuf_1 \gen_obs_vmem[128].sdcbuf_gen_vmem  (.A(\vmem[128] ),
    .X(\vmem_after_buf[128] ));
 clkbuf_1 \gen_obs_vmem[129].sdcbuf_gen_vmem  (.A(\vmem[129] ),
    .X(\vmem_after_buf[129] ));
 clkbuf_1 \gen_obs_vmem[12].sdcbuf_gen_vmem  (.A(\vmem[12] ),
    .X(\vmem_after_buf[12] ));
 clkbuf_1 \gen_obs_vmem[130].sdcbuf_gen_vmem  (.A(\vmem[130] ),
    .X(\vmem_after_buf[130] ));
 clkbuf_1 \gen_obs_vmem[131].sdcbuf_gen_vmem  (.A(\vmem[131] ),
    .X(\vmem_after_buf[131] ));
 clkbuf_1 \gen_obs_vmem[132].sdcbuf_gen_vmem  (.A(\vmem[132] ),
    .X(\vmem_after_buf[132] ));
 clkbuf_1 \gen_obs_vmem[133].sdcbuf_gen_vmem  (.A(\vmem[133] ),
    .X(\vmem_after_buf[133] ));
 clkbuf_1 \gen_obs_vmem[134].sdcbuf_gen_vmem  (.A(\vmem[134] ),
    .X(\vmem_after_buf[134] ));
 clkbuf_1 \gen_obs_vmem[135].sdcbuf_gen_vmem  (.A(\vmem[135] ),
    .X(\vmem_after_buf[135] ));
 clkbuf_1 \gen_obs_vmem[136].sdcbuf_gen_vmem  (.A(\vmem[136] ),
    .X(\vmem_after_buf[136] ));
 clkbuf_1 \gen_obs_vmem[137].sdcbuf_gen_vmem  (.A(\vmem[137] ),
    .X(\vmem_after_buf[137] ));
 clkbuf_1 \gen_obs_vmem[138].sdcbuf_gen_vmem  (.A(\vmem[138] ),
    .X(\vmem_after_buf[138] ));
 clkbuf_1 \gen_obs_vmem[139].sdcbuf_gen_vmem  (.A(\vmem[139] ),
    .X(\vmem_after_buf[139] ));
 clkbuf_1 \gen_obs_vmem[13].sdcbuf_gen_vmem  (.A(\vmem[13] ),
    .X(\vmem_after_buf[13] ));
 clkbuf_1 \gen_obs_vmem[140].sdcbuf_gen_vmem  (.A(\vmem[140] ),
    .X(\vmem_after_buf[140] ));
 clkbuf_1 \gen_obs_vmem[141].sdcbuf_gen_vmem  (.A(\vmem[141] ),
    .X(\vmem_after_buf[141] ));
 clkbuf_1 \gen_obs_vmem[142].sdcbuf_gen_vmem  (.A(\vmem[142] ),
    .X(\vmem_after_buf[142] ));
 clkbuf_1 \gen_obs_vmem[143].sdcbuf_gen_vmem  (.A(\vmem[143] ),
    .X(\vmem_after_buf[143] ));
 clkbuf_1 \gen_obs_vmem[144].sdcbuf_gen_vmem  (.A(\vmem[144] ),
    .X(\vmem_after_buf[144] ));
 clkbuf_1 \gen_obs_vmem[145].sdcbuf_gen_vmem  (.A(\vmem[145] ),
    .X(\vmem_after_buf[145] ));
 clkbuf_1 \gen_obs_vmem[146].sdcbuf_gen_vmem  (.A(\vmem[146] ),
    .X(\vmem_after_buf[146] ));
 clkbuf_1 \gen_obs_vmem[147].sdcbuf_gen_vmem  (.A(\vmem[147] ),
    .X(\vmem_after_buf[147] ));
 clkbuf_1 \gen_obs_vmem[148].sdcbuf_gen_vmem  (.A(\vmem[148] ),
    .X(\vmem_after_buf[148] ));
 clkbuf_1 \gen_obs_vmem[149].sdcbuf_gen_vmem  (.A(\vmem[149] ),
    .X(\vmem_after_buf[149] ));
 clkbuf_1 \gen_obs_vmem[14].sdcbuf_gen_vmem  (.A(\vmem[14] ),
    .X(\vmem_after_buf[14] ));
 clkbuf_1 \gen_obs_vmem[150].sdcbuf_gen_vmem  (.A(\vmem[150] ),
    .X(\vmem_after_buf[150] ));
 clkbuf_1 \gen_obs_vmem[151].sdcbuf_gen_vmem  (.A(\vmem[151] ),
    .X(\vmem_after_buf[151] ));
 clkbuf_1 \gen_obs_vmem[152].sdcbuf_gen_vmem  (.A(\vmem[152] ),
    .X(\vmem_after_buf[152] ));
 clkbuf_1 \gen_obs_vmem[153].sdcbuf_gen_vmem  (.A(\vmem[153] ),
    .X(\vmem_after_buf[153] ));
 clkbuf_1 \gen_obs_vmem[154].sdcbuf_gen_vmem  (.A(\vmem[154] ),
    .X(\vmem_after_buf[154] ));
 clkbuf_1 \gen_obs_vmem[155].sdcbuf_gen_vmem  (.A(\vmem[155] ),
    .X(\vmem_after_buf[155] ));
 clkbuf_1 \gen_obs_vmem[156].sdcbuf_gen_vmem  (.A(\vmem[156] ),
    .X(\vmem_after_buf[156] ));
 clkbuf_1 \gen_obs_vmem[157].sdcbuf_gen_vmem  (.A(\vmem[157] ),
    .X(\vmem_after_buf[157] ));
 clkbuf_1 \gen_obs_vmem[158].sdcbuf_gen_vmem  (.A(\vmem[158] ),
    .X(\vmem_after_buf[158] ));
 clkbuf_1 \gen_obs_vmem[159].sdcbuf_gen_vmem  (.A(\vmem[159] ),
    .X(\vmem_after_buf[159] ));
 clkbuf_1 \gen_obs_vmem[15].sdcbuf_gen_vmem  (.A(\vmem[15] ),
    .X(\vmem_after_buf[15] ));
 clkbuf_1 \gen_obs_vmem[160].sdcbuf_gen_vmem  (.A(\vmem[160] ),
    .X(\vmem_after_buf[160] ));
 clkbuf_1 \gen_obs_vmem[161].sdcbuf_gen_vmem  (.A(\vmem[161] ),
    .X(\vmem_after_buf[161] ));
 clkbuf_1 \gen_obs_vmem[162].sdcbuf_gen_vmem  (.A(\vmem[162] ),
    .X(\vmem_after_buf[162] ));
 clkbuf_1 \gen_obs_vmem[163].sdcbuf_gen_vmem  (.A(\vmem[163] ),
    .X(\vmem_after_buf[163] ));
 clkbuf_1 \gen_obs_vmem[164].sdcbuf_gen_vmem  (.A(\vmem[164] ),
    .X(\vmem_after_buf[164] ));
 clkbuf_1 \gen_obs_vmem[165].sdcbuf_gen_vmem  (.A(\vmem[165] ),
    .X(\vmem_after_buf[165] ));
 clkbuf_1 \gen_obs_vmem[166].sdcbuf_gen_vmem  (.A(\vmem[166] ),
    .X(\vmem_after_buf[166] ));
 clkbuf_1 \gen_obs_vmem[167].sdcbuf_gen_vmem  (.A(\vmem[167] ),
    .X(\vmem_after_buf[167] ));
 clkbuf_1 \gen_obs_vmem[168].sdcbuf_gen_vmem  (.A(\vmem[168] ),
    .X(\vmem_after_buf[168] ));
 clkbuf_1 \gen_obs_vmem[169].sdcbuf_gen_vmem  (.A(\vmem[169] ),
    .X(\vmem_after_buf[169] ));
 clkbuf_1 \gen_obs_vmem[16].sdcbuf_gen_vmem  (.A(\vmem[16] ),
    .X(\vmem_after_buf[16] ));
 clkbuf_1 \gen_obs_vmem[170].sdcbuf_gen_vmem  (.A(\vmem[170] ),
    .X(\vmem_after_buf[170] ));
 clkbuf_1 \gen_obs_vmem[171].sdcbuf_gen_vmem  (.A(\vmem[171] ),
    .X(\vmem_after_buf[171] ));
 clkbuf_1 \gen_obs_vmem[172].sdcbuf_gen_vmem  (.A(\vmem[172] ),
    .X(\vmem_after_buf[172] ));
 clkbuf_1 \gen_obs_vmem[173].sdcbuf_gen_vmem  (.A(\vmem[173] ),
    .X(\vmem_after_buf[173] ));
 clkbuf_1 \gen_obs_vmem[174].sdcbuf_gen_vmem  (.A(\vmem[174] ),
    .X(\vmem_after_buf[174] ));
 clkbuf_1 \gen_obs_vmem[175].sdcbuf_gen_vmem  (.A(\vmem[175] ),
    .X(\vmem_after_buf[175] ));
 clkbuf_1 \gen_obs_vmem[176].sdcbuf_gen_vmem  (.A(\vmem[176] ),
    .X(\vmem_after_buf[176] ));
 clkbuf_1 \gen_obs_vmem[177].sdcbuf_gen_vmem  (.A(\vmem[177] ),
    .X(\vmem_after_buf[177] ));
 clkbuf_1 \gen_obs_vmem[178].sdcbuf_gen_vmem  (.A(\vmem[178] ),
    .X(\vmem_after_buf[178] ));
 clkbuf_1 \gen_obs_vmem[179].sdcbuf_gen_vmem  (.A(\vmem[179] ),
    .X(\vmem_after_buf[179] ));
 clkbuf_1 \gen_obs_vmem[17].sdcbuf_gen_vmem  (.A(\vmem[17] ),
    .X(\vmem_after_buf[17] ));
 clkbuf_1 \gen_obs_vmem[180].sdcbuf_gen_vmem  (.A(\vmem[180] ),
    .X(\vmem_after_buf[180] ));
 clkbuf_1 \gen_obs_vmem[181].sdcbuf_gen_vmem  (.A(\vmem[181] ),
    .X(\vmem_after_buf[181] ));
 clkbuf_1 \gen_obs_vmem[182].sdcbuf_gen_vmem  (.A(\vmem[182] ),
    .X(\vmem_after_buf[182] ));
 clkbuf_1 \gen_obs_vmem[183].sdcbuf_gen_vmem  (.A(\vmem[183] ),
    .X(\vmem_after_buf[183] ));
 clkbuf_1 \gen_obs_vmem[184].sdcbuf_gen_vmem  (.A(\vmem[184] ),
    .X(\vmem_after_buf[184] ));
 clkbuf_1 \gen_obs_vmem[185].sdcbuf_gen_vmem  (.A(\vmem[185] ),
    .X(\vmem_after_buf[185] ));
 clkbuf_1 \gen_obs_vmem[186].sdcbuf_gen_vmem  (.A(\vmem[186] ),
    .X(\vmem_after_buf[186] ));
 clkbuf_1 \gen_obs_vmem[187].sdcbuf_gen_vmem  (.A(\vmem[187] ),
    .X(\vmem_after_buf[187] ));
 clkbuf_1 \gen_obs_vmem[188].sdcbuf_gen_vmem  (.A(\vmem[188] ),
    .X(\vmem_after_buf[188] ));
 clkbuf_1 \gen_obs_vmem[189].sdcbuf_gen_vmem  (.A(\vmem[189] ),
    .X(\vmem_after_buf[189] ));
 clkbuf_1 \gen_obs_vmem[18].sdcbuf_gen_vmem  (.A(\vmem[18] ),
    .X(\vmem_after_buf[18] ));
 clkbuf_1 \gen_obs_vmem[190].sdcbuf_gen_vmem  (.A(\vmem[190] ),
    .X(\vmem_after_buf[190] ));
 clkbuf_1 \gen_obs_vmem[191].sdcbuf_gen_vmem  (.A(\vmem[191] ),
    .X(\vmem_after_buf[191] ));
 clkbuf_1 \gen_obs_vmem[192].sdcbuf_gen_vmem  (.A(\vmem[192] ),
    .X(\vmem_after_buf[192] ));
 clkbuf_1 \gen_obs_vmem[193].sdcbuf_gen_vmem  (.A(\vmem[193] ),
    .X(\vmem_after_buf[193] ));
 clkbuf_1 \gen_obs_vmem[194].sdcbuf_gen_vmem  (.A(\vmem[194] ),
    .X(\vmem_after_buf[194] ));
 clkbuf_1 \gen_obs_vmem[195].sdcbuf_gen_vmem  (.A(\vmem[195] ),
    .X(\vmem_after_buf[195] ));
 clkbuf_1 \gen_obs_vmem[196].sdcbuf_gen_vmem  (.A(\vmem[196] ),
    .X(\vmem_after_buf[196] ));
 clkbuf_1 \gen_obs_vmem[197].sdcbuf_gen_vmem  (.A(\vmem[197] ),
    .X(\vmem_after_buf[197] ));
 clkbuf_1 \gen_obs_vmem[198].sdcbuf_gen_vmem  (.A(\vmem[198] ),
    .X(\vmem_after_buf[198] ));
 clkbuf_1 \gen_obs_vmem[199].sdcbuf_gen_vmem  (.A(\vmem[199] ),
    .X(\vmem_after_buf[199] ));
 clkbuf_1 \gen_obs_vmem[19].sdcbuf_gen_vmem  (.A(\vmem[19] ),
    .X(\vmem_after_buf[19] ));
 clkbuf_1 \gen_obs_vmem[1].sdcbuf_gen_vmem  (.A(\vmem[1] ),
    .X(\vmem_after_buf[1] ));
 clkbuf_1 \gen_obs_vmem[200].sdcbuf_gen_vmem  (.A(\vmem[200] ),
    .X(\vmem_after_buf[200] ));
 clkbuf_1 \gen_obs_vmem[201].sdcbuf_gen_vmem  (.A(\vmem[201] ),
    .X(\vmem_after_buf[201] ));
 clkbuf_1 \gen_obs_vmem[202].sdcbuf_gen_vmem  (.A(\vmem[202] ),
    .X(\vmem_after_buf[202] ));
 clkbuf_1 \gen_obs_vmem[203].sdcbuf_gen_vmem  (.A(\vmem[203] ),
    .X(\vmem_after_buf[203] ));
 clkbuf_1 \gen_obs_vmem[204].sdcbuf_gen_vmem  (.A(\vmem[204] ),
    .X(\vmem_after_buf[204] ));
 clkbuf_1 \gen_obs_vmem[205].sdcbuf_gen_vmem  (.A(\vmem[205] ),
    .X(\vmem_after_buf[205] ));
 clkbuf_1 \gen_obs_vmem[206].sdcbuf_gen_vmem  (.A(\vmem[206] ),
    .X(\vmem_after_buf[206] ));
 clkbuf_1 \gen_obs_vmem[207].sdcbuf_gen_vmem  (.A(\vmem[207] ),
    .X(\vmem_after_buf[207] ));
 clkbuf_1 \gen_obs_vmem[208].sdcbuf_gen_vmem  (.A(\vmem[208] ),
    .X(\vmem_after_buf[208] ));
 clkbuf_1 \gen_obs_vmem[209].sdcbuf_gen_vmem  (.A(\vmem[209] ),
    .X(\vmem_after_buf[209] ));
 clkbuf_1 \gen_obs_vmem[20].sdcbuf_gen_vmem  (.A(\vmem[20] ),
    .X(\vmem_after_buf[20] ));
 clkbuf_1 \gen_obs_vmem[210].sdcbuf_gen_vmem  (.A(\vmem[210] ),
    .X(\vmem_after_buf[210] ));
 clkbuf_1 \gen_obs_vmem[211].sdcbuf_gen_vmem  (.A(\vmem[211] ),
    .X(\vmem_after_buf[211] ));
 clkbuf_1 \gen_obs_vmem[212].sdcbuf_gen_vmem  (.A(\vmem[212] ),
    .X(\vmem_after_buf[212] ));
 clkbuf_1 \gen_obs_vmem[213].sdcbuf_gen_vmem  (.A(\vmem[213] ),
    .X(\vmem_after_buf[213] ));
 clkbuf_1 \gen_obs_vmem[214].sdcbuf_gen_vmem  (.A(\vmem[214] ),
    .X(\vmem_after_buf[214] ));
 clkbuf_1 \gen_obs_vmem[215].sdcbuf_gen_vmem  (.A(\vmem[215] ),
    .X(\vmem_after_buf[215] ));
 clkbuf_1 \gen_obs_vmem[216].sdcbuf_gen_vmem  (.A(\vmem[216] ),
    .X(\vmem_after_buf[216] ));
 clkbuf_1 \gen_obs_vmem[217].sdcbuf_gen_vmem  (.A(\vmem[217] ),
    .X(\vmem_after_buf[217] ));
 clkbuf_1 \gen_obs_vmem[218].sdcbuf_gen_vmem  (.A(\vmem[218] ),
    .X(\vmem_after_buf[218] ));
 clkbuf_1 \gen_obs_vmem[219].sdcbuf_gen_vmem  (.A(\vmem[219] ),
    .X(\vmem_after_buf[219] ));
 clkbuf_1 \gen_obs_vmem[21].sdcbuf_gen_vmem  (.A(\vmem[21] ),
    .X(\vmem_after_buf[21] ));
 clkbuf_1 \gen_obs_vmem[220].sdcbuf_gen_vmem  (.A(\vmem[220] ),
    .X(\vmem_after_buf[220] ));
 clkbuf_1 \gen_obs_vmem[221].sdcbuf_gen_vmem  (.A(\vmem[221] ),
    .X(\vmem_after_buf[221] ));
 clkbuf_1 \gen_obs_vmem[222].sdcbuf_gen_vmem  (.A(\vmem[222] ),
    .X(\vmem_after_buf[222] ));
 clkbuf_1 \gen_obs_vmem[223].sdcbuf_gen_vmem  (.A(\vmem[223] ),
    .X(\vmem_after_buf[223] ));
 clkbuf_1 \gen_obs_vmem[224].sdcbuf_gen_vmem  (.A(\vmem[224] ),
    .X(\vmem_after_buf[224] ));
 clkbuf_1 \gen_obs_vmem[225].sdcbuf_gen_vmem  (.A(\vmem[225] ),
    .X(\vmem_after_buf[225] ));
 clkbuf_1 \gen_obs_vmem[226].sdcbuf_gen_vmem  (.A(\vmem[226] ),
    .X(\vmem_after_buf[226] ));
 clkbuf_1 \gen_obs_vmem[227].sdcbuf_gen_vmem  (.A(\vmem[227] ),
    .X(\vmem_after_buf[227] ));
 clkbuf_1 \gen_obs_vmem[228].sdcbuf_gen_vmem  (.A(\vmem[228] ),
    .X(\vmem_after_buf[228] ));
 clkbuf_1 \gen_obs_vmem[229].sdcbuf_gen_vmem  (.A(\vmem[229] ),
    .X(\vmem_after_buf[229] ));
 clkbuf_1 \gen_obs_vmem[22].sdcbuf_gen_vmem  (.A(\vmem[22] ),
    .X(\vmem_after_buf[22] ));
 clkbuf_1 \gen_obs_vmem[230].sdcbuf_gen_vmem  (.A(\vmem[230] ),
    .X(\vmem_after_buf[230] ));
 clkbuf_1 \gen_obs_vmem[231].sdcbuf_gen_vmem  (.A(\vmem[231] ),
    .X(\vmem_after_buf[231] ));
 clkbuf_1 \gen_obs_vmem[232].sdcbuf_gen_vmem  (.A(\vmem[232] ),
    .X(\vmem_after_buf[232] ));
 clkbuf_1 \gen_obs_vmem[233].sdcbuf_gen_vmem  (.A(\vmem[233] ),
    .X(\vmem_after_buf[233] ));
 clkbuf_1 \gen_obs_vmem[234].sdcbuf_gen_vmem  (.A(\vmem[234] ),
    .X(\vmem_after_buf[234] ));
 clkbuf_1 \gen_obs_vmem[235].sdcbuf_gen_vmem  (.A(\vmem[235] ),
    .X(\vmem_after_buf[235] ));
 clkbuf_1 \gen_obs_vmem[236].sdcbuf_gen_vmem  (.A(\vmem[236] ),
    .X(\vmem_after_buf[236] ));
 clkbuf_1 \gen_obs_vmem[237].sdcbuf_gen_vmem  (.A(\vmem[237] ),
    .X(\vmem_after_buf[237] ));
 clkbuf_1 \gen_obs_vmem[238].sdcbuf_gen_vmem  (.A(\vmem[238] ),
    .X(\vmem_after_buf[238] ));
 clkbuf_1 \gen_obs_vmem[239].sdcbuf_gen_vmem  (.A(\vmem[239] ),
    .X(\vmem_after_buf[239] ));
 clkbuf_1 \gen_obs_vmem[23].sdcbuf_gen_vmem  (.A(\vmem[23] ),
    .X(\vmem_after_buf[23] ));
 clkbuf_1 \gen_obs_vmem[240].sdcbuf_gen_vmem  (.A(\vmem[240] ),
    .X(\vmem_after_buf[240] ));
 clkbuf_1 \gen_obs_vmem[241].sdcbuf_gen_vmem  (.A(\vmem[241] ),
    .X(\vmem_after_buf[241] ));
 clkbuf_1 \gen_obs_vmem[242].sdcbuf_gen_vmem  (.A(\vmem[242] ),
    .X(\vmem_after_buf[242] ));
 clkbuf_1 \gen_obs_vmem[243].sdcbuf_gen_vmem  (.A(\vmem[243] ),
    .X(\vmem_after_buf[243] ));
 clkbuf_1 \gen_obs_vmem[244].sdcbuf_gen_vmem  (.A(\vmem[244] ),
    .X(\vmem_after_buf[244] ));
 clkbuf_1 \gen_obs_vmem[245].sdcbuf_gen_vmem  (.A(\vmem[245] ),
    .X(\vmem_after_buf[245] ));
 clkbuf_1 \gen_obs_vmem[246].sdcbuf_gen_vmem  (.A(\vmem[246] ),
    .X(\vmem_after_buf[246] ));
 clkbuf_1 \gen_obs_vmem[247].sdcbuf_gen_vmem  (.A(\vmem[247] ),
    .X(\vmem_after_buf[247] ));
 clkbuf_1 \gen_obs_vmem[248].sdcbuf_gen_vmem  (.A(\vmem[248] ),
    .X(\vmem_after_buf[248] ));
 clkbuf_1 \gen_obs_vmem[249].sdcbuf_gen_vmem  (.A(\vmem[249] ),
    .X(\vmem_after_buf[249] ));
 clkbuf_1 \gen_obs_vmem[24].sdcbuf_gen_vmem  (.A(\vmem[24] ),
    .X(\vmem_after_buf[24] ));
 clkbuf_1 \gen_obs_vmem[250].sdcbuf_gen_vmem  (.A(\vmem[250] ),
    .X(\vmem_after_buf[250] ));
 clkbuf_1 \gen_obs_vmem[251].sdcbuf_gen_vmem  (.A(\vmem[251] ),
    .X(\vmem_after_buf[251] ));
 clkbuf_1 \gen_obs_vmem[252].sdcbuf_gen_vmem  (.A(\vmem[252] ),
    .X(\vmem_after_buf[252] ));
 clkbuf_1 \gen_obs_vmem[253].sdcbuf_gen_vmem  (.A(\vmem[253] ),
    .X(\vmem_after_buf[253] ));
 clkbuf_1 \gen_obs_vmem[254].sdcbuf_gen_vmem  (.A(\vmem[254] ),
    .X(\vmem_after_buf[254] ));
 clkbuf_1 \gen_obs_vmem[255].sdcbuf_gen_vmem  (.A(\vmem[255] ),
    .X(\vmem_after_buf[255] ));
 clkbuf_1 \gen_obs_vmem[256].sdcbuf_gen_vmem  (.A(\vmem[256] ),
    .X(\vmem_after_buf[256] ));
 clkbuf_1 \gen_obs_vmem[257].sdcbuf_gen_vmem  (.A(\vmem[257] ),
    .X(\vmem_after_buf[257] ));
 clkbuf_1 \gen_obs_vmem[258].sdcbuf_gen_vmem  (.A(\vmem[258] ),
    .X(\vmem_after_buf[258] ));
 clkbuf_1 \gen_obs_vmem[259].sdcbuf_gen_vmem  (.A(\vmem[259] ),
    .X(\vmem_after_buf[259] ));
 clkbuf_1 \gen_obs_vmem[25].sdcbuf_gen_vmem  (.A(\vmem[25] ),
    .X(\vmem_after_buf[25] ));
 clkbuf_1 \gen_obs_vmem[260].sdcbuf_gen_vmem  (.A(\vmem[260] ),
    .X(\vmem_after_buf[260] ));
 clkbuf_1 \gen_obs_vmem[261].sdcbuf_gen_vmem  (.A(\vmem[261] ),
    .X(\vmem_after_buf[261] ));
 clkbuf_1 \gen_obs_vmem[262].sdcbuf_gen_vmem  (.A(\vmem[262] ),
    .X(\vmem_after_buf[262] ));
 clkbuf_1 \gen_obs_vmem[263].sdcbuf_gen_vmem  (.A(\vmem[263] ),
    .X(\vmem_after_buf[263] ));
 clkbuf_1 \gen_obs_vmem[264].sdcbuf_gen_vmem  (.A(\vmem[264] ),
    .X(\vmem_after_buf[264] ));
 clkbuf_1 \gen_obs_vmem[265].sdcbuf_gen_vmem  (.A(\vmem[265] ),
    .X(\vmem_after_buf[265] ));
 clkbuf_1 \gen_obs_vmem[266].sdcbuf_gen_vmem  (.A(\vmem[266] ),
    .X(\vmem_after_buf[266] ));
 clkbuf_1 \gen_obs_vmem[267].sdcbuf_gen_vmem  (.A(\vmem[267] ),
    .X(\vmem_after_buf[267] ));
 clkbuf_1 \gen_obs_vmem[268].sdcbuf_gen_vmem  (.A(\vmem[268] ),
    .X(\vmem_after_buf[268] ));
 clkbuf_1 \gen_obs_vmem[269].sdcbuf_gen_vmem  (.A(\vmem[269] ),
    .X(\vmem_after_buf[269] ));
 clkbuf_1 \gen_obs_vmem[26].sdcbuf_gen_vmem  (.A(\vmem[26] ),
    .X(\vmem_after_buf[26] ));
 clkbuf_1 \gen_obs_vmem[270].sdcbuf_gen_vmem  (.A(\vmem[270] ),
    .X(\vmem_after_buf[270] ));
 clkbuf_1 \gen_obs_vmem[271].sdcbuf_gen_vmem  (.A(\vmem[271] ),
    .X(\vmem_after_buf[271] ));
 clkbuf_1 \gen_obs_vmem[272].sdcbuf_gen_vmem  (.A(\vmem[272] ),
    .X(\vmem_after_buf[272] ));
 clkbuf_1 \gen_obs_vmem[273].sdcbuf_gen_vmem  (.A(\vmem[273] ),
    .X(\vmem_after_buf[273] ));
 clkbuf_1 \gen_obs_vmem[274].sdcbuf_gen_vmem  (.A(\vmem[274] ),
    .X(\vmem_after_buf[274] ));
 clkbuf_1 \gen_obs_vmem[275].sdcbuf_gen_vmem  (.A(\vmem[275] ),
    .X(\vmem_after_buf[275] ));
 clkbuf_1 \gen_obs_vmem[276].sdcbuf_gen_vmem  (.A(\vmem[276] ),
    .X(\vmem_after_buf[276] ));
 clkbuf_1 \gen_obs_vmem[277].sdcbuf_gen_vmem  (.A(\vmem[277] ),
    .X(\vmem_after_buf[277] ));
 clkbuf_1 \gen_obs_vmem[278].sdcbuf_gen_vmem  (.A(\vmem[278] ),
    .X(\vmem_after_buf[278] ));
 clkbuf_1 \gen_obs_vmem[279].sdcbuf_gen_vmem  (.A(\vmem[279] ),
    .X(\vmem_after_buf[279] ));
 clkbuf_1 \gen_obs_vmem[27].sdcbuf_gen_vmem  (.A(\vmem[27] ),
    .X(\vmem_after_buf[27] ));
 clkbuf_1 \gen_obs_vmem[280].sdcbuf_gen_vmem  (.A(\vmem[280] ),
    .X(\vmem_after_buf[280] ));
 clkbuf_1 \gen_obs_vmem[281].sdcbuf_gen_vmem  (.A(\vmem[281] ),
    .X(\vmem_after_buf[281] ));
 clkbuf_1 \gen_obs_vmem[282].sdcbuf_gen_vmem  (.A(\vmem[282] ),
    .X(\vmem_after_buf[282] ));
 clkbuf_1 \gen_obs_vmem[283].sdcbuf_gen_vmem  (.A(\vmem[283] ),
    .X(\vmem_after_buf[283] ));
 clkbuf_1 \gen_obs_vmem[284].sdcbuf_gen_vmem  (.A(\vmem[284] ),
    .X(\vmem_after_buf[284] ));
 clkbuf_1 \gen_obs_vmem[285].sdcbuf_gen_vmem  (.A(\vmem[285] ),
    .X(\vmem_after_buf[285] ));
 clkbuf_1 \gen_obs_vmem[286].sdcbuf_gen_vmem  (.A(\vmem[286] ),
    .X(\vmem_after_buf[286] ));
 clkbuf_1 \gen_obs_vmem[287].sdcbuf_gen_vmem  (.A(\vmem[287] ),
    .X(\vmem_after_buf[287] ));
 clkbuf_1 \gen_obs_vmem[288].sdcbuf_gen_vmem  (.A(\vmem[288] ),
    .X(\vmem_after_buf[288] ));
 clkbuf_1 \gen_obs_vmem[289].sdcbuf_gen_vmem  (.A(\vmem[289] ),
    .X(\vmem_after_buf[289] ));
 clkbuf_1 \gen_obs_vmem[28].sdcbuf_gen_vmem  (.A(\vmem[28] ),
    .X(\vmem_after_buf[28] ));
 clkbuf_1 \gen_obs_vmem[290].sdcbuf_gen_vmem  (.A(\vmem[290] ),
    .X(\vmem_after_buf[290] ));
 clkbuf_1 \gen_obs_vmem[291].sdcbuf_gen_vmem  (.A(\vmem[291] ),
    .X(\vmem_after_buf[291] ));
 clkbuf_1 \gen_obs_vmem[292].sdcbuf_gen_vmem  (.A(\vmem[292] ),
    .X(\vmem_after_buf[292] ));
 clkbuf_1 \gen_obs_vmem[293].sdcbuf_gen_vmem  (.A(\vmem[293] ),
    .X(\vmem_after_buf[293] ));
 clkbuf_1 \gen_obs_vmem[294].sdcbuf_gen_vmem  (.A(\vmem[294] ),
    .X(\vmem_after_buf[294] ));
 clkbuf_1 \gen_obs_vmem[295].sdcbuf_gen_vmem  (.A(\vmem[295] ),
    .X(\vmem_after_buf[295] ));
 clkbuf_1 \gen_obs_vmem[296].sdcbuf_gen_vmem  (.A(\vmem[296] ),
    .X(\vmem_after_buf[296] ));
 clkbuf_1 \gen_obs_vmem[297].sdcbuf_gen_vmem  (.A(\vmem[297] ),
    .X(\vmem_after_buf[297] ));
 clkbuf_1 \gen_obs_vmem[298].sdcbuf_gen_vmem  (.A(\vmem[298] ),
    .X(\vmem_after_buf[298] ));
 clkbuf_1 \gen_obs_vmem[299].sdcbuf_gen_vmem  (.A(\vmem[299] ),
    .X(\vmem_after_buf[299] ));
 clkbuf_1 \gen_obs_vmem[29].sdcbuf_gen_vmem  (.A(\vmem[29] ),
    .X(\vmem_after_buf[29] ));
 clkbuf_1 \gen_obs_vmem[2].sdcbuf_gen_vmem  (.A(\vmem[2] ),
    .X(\vmem_after_buf[2] ));
 clkbuf_1 \gen_obs_vmem[300].sdcbuf_gen_vmem  (.A(\vmem[300] ),
    .X(\vmem_after_buf[300] ));
 clkbuf_1 \gen_obs_vmem[301].sdcbuf_gen_vmem  (.A(\vmem[301] ),
    .X(\vmem_after_buf[301] ));
 clkbuf_1 \gen_obs_vmem[302].sdcbuf_gen_vmem  (.A(\vmem[302] ),
    .X(\vmem_after_buf[302] ));
 clkbuf_1 \gen_obs_vmem[303].sdcbuf_gen_vmem  (.A(\vmem[303] ),
    .X(\vmem_after_buf[303] ));
 clkbuf_1 \gen_obs_vmem[304].sdcbuf_gen_vmem  (.A(\vmem[304] ),
    .X(\vmem_after_buf[304] ));
 clkbuf_1 \gen_obs_vmem[305].sdcbuf_gen_vmem  (.A(\vmem[305] ),
    .X(\vmem_after_buf[305] ));
 clkbuf_1 \gen_obs_vmem[306].sdcbuf_gen_vmem  (.A(\vmem[306] ),
    .X(\vmem_after_buf[306] ));
 clkbuf_1 \gen_obs_vmem[307].sdcbuf_gen_vmem  (.A(\vmem[307] ),
    .X(\vmem_after_buf[307] ));
 clkbuf_1 \gen_obs_vmem[308].sdcbuf_gen_vmem  (.A(\vmem[308] ),
    .X(\vmem_after_buf[308] ));
 clkbuf_1 \gen_obs_vmem[309].sdcbuf_gen_vmem  (.A(\vmem[309] ),
    .X(\vmem_after_buf[309] ));
 clkbuf_1 \gen_obs_vmem[30].sdcbuf_gen_vmem  (.A(\vmem[30] ),
    .X(\vmem_after_buf[30] ));
 clkbuf_1 \gen_obs_vmem[310].sdcbuf_gen_vmem  (.A(\vmem[310] ),
    .X(\vmem_after_buf[310] ));
 clkbuf_1 \gen_obs_vmem[311].sdcbuf_gen_vmem  (.A(\vmem[311] ),
    .X(\vmem_after_buf[311] ));
 clkbuf_1 \gen_obs_vmem[312].sdcbuf_gen_vmem  (.A(\vmem[312] ),
    .X(\vmem_after_buf[312] ));
 clkbuf_1 \gen_obs_vmem[313].sdcbuf_gen_vmem  (.A(\vmem[313] ),
    .X(\vmem_after_buf[313] ));
 clkbuf_1 \gen_obs_vmem[314].sdcbuf_gen_vmem  (.A(\vmem[314] ),
    .X(\vmem_after_buf[314] ));
 clkbuf_1 \gen_obs_vmem[315].sdcbuf_gen_vmem  (.A(\vmem[315] ),
    .X(\vmem_after_buf[315] ));
 clkbuf_1 \gen_obs_vmem[316].sdcbuf_gen_vmem  (.A(\vmem[316] ),
    .X(\vmem_after_buf[316] ));
 clkbuf_1 \gen_obs_vmem[317].sdcbuf_gen_vmem  (.A(\vmem[317] ),
    .X(\vmem_after_buf[317] ));
 clkbuf_1 \gen_obs_vmem[318].sdcbuf_gen_vmem  (.A(\vmem[318] ),
    .X(\vmem_after_buf[318] ));
 clkbuf_1 \gen_obs_vmem[319].sdcbuf_gen_vmem  (.A(\vmem[319] ),
    .X(\vmem_after_buf[319] ));
 clkbuf_1 \gen_obs_vmem[31].sdcbuf_gen_vmem  (.A(\vmem[31] ),
    .X(\vmem_after_buf[31] ));
 clkbuf_1 \gen_obs_vmem[320].sdcbuf_gen_vmem  (.A(\vmem[320] ),
    .X(\vmem_after_buf[320] ));
 clkbuf_1 \gen_obs_vmem[321].sdcbuf_gen_vmem  (.A(\vmem[321] ),
    .X(\vmem_after_buf[321] ));
 clkbuf_1 \gen_obs_vmem[322].sdcbuf_gen_vmem  (.A(\vmem[322] ),
    .X(\vmem_after_buf[322] ));
 clkbuf_1 \gen_obs_vmem[323].sdcbuf_gen_vmem  (.A(\vmem[323] ),
    .X(\vmem_after_buf[323] ));
 clkbuf_1 \gen_obs_vmem[324].sdcbuf_gen_vmem  (.A(\vmem[324] ),
    .X(\vmem_after_buf[324] ));
 clkbuf_1 \gen_obs_vmem[325].sdcbuf_gen_vmem  (.A(\vmem[325] ),
    .X(\vmem_after_buf[325] ));
 clkbuf_1 \gen_obs_vmem[326].sdcbuf_gen_vmem  (.A(\vmem[326] ),
    .X(\vmem_after_buf[326] ));
 clkbuf_1 \gen_obs_vmem[327].sdcbuf_gen_vmem  (.A(\vmem[327] ),
    .X(\vmem_after_buf[327] ));
 clkbuf_1 \gen_obs_vmem[328].sdcbuf_gen_vmem  (.A(\vmem[328] ),
    .X(\vmem_after_buf[328] ));
 clkbuf_1 \gen_obs_vmem[329].sdcbuf_gen_vmem  (.A(\vmem[329] ),
    .X(\vmem_after_buf[329] ));
 clkbuf_1 \gen_obs_vmem[32].sdcbuf_gen_vmem  (.A(\vmem[32] ),
    .X(\vmem_after_buf[32] ));
 clkbuf_1 \gen_obs_vmem[330].sdcbuf_gen_vmem  (.A(\vmem[330] ),
    .X(\vmem_after_buf[330] ));
 clkbuf_1 \gen_obs_vmem[331].sdcbuf_gen_vmem  (.A(\vmem[331] ),
    .X(\vmem_after_buf[331] ));
 clkbuf_1 \gen_obs_vmem[332].sdcbuf_gen_vmem  (.A(\vmem[332] ),
    .X(\vmem_after_buf[332] ));
 clkbuf_1 \gen_obs_vmem[333].sdcbuf_gen_vmem  (.A(\vmem[333] ),
    .X(\vmem_after_buf[333] ));
 clkbuf_1 \gen_obs_vmem[334].sdcbuf_gen_vmem  (.A(\vmem[334] ),
    .X(\vmem_after_buf[334] ));
 clkbuf_1 \gen_obs_vmem[335].sdcbuf_gen_vmem  (.A(\vmem[335] ),
    .X(\vmem_after_buf[335] ));
 clkbuf_1 \gen_obs_vmem[336].sdcbuf_gen_vmem  (.A(\vmem[336] ),
    .X(\vmem_after_buf[336] ));
 clkbuf_1 \gen_obs_vmem[337].sdcbuf_gen_vmem  (.A(\vmem[337] ),
    .X(\vmem_after_buf[337] ));
 clkbuf_1 \gen_obs_vmem[338].sdcbuf_gen_vmem  (.A(\vmem[338] ),
    .X(\vmem_after_buf[338] ));
 clkbuf_1 \gen_obs_vmem[339].sdcbuf_gen_vmem  (.A(\vmem[339] ),
    .X(\vmem_after_buf[339] ));
 clkbuf_1 \gen_obs_vmem[33].sdcbuf_gen_vmem  (.A(\vmem[33] ),
    .X(\vmem_after_buf[33] ));
 clkbuf_1 \gen_obs_vmem[340].sdcbuf_gen_vmem  (.A(\vmem[340] ),
    .X(\vmem_after_buf[340] ));
 clkbuf_1 \gen_obs_vmem[341].sdcbuf_gen_vmem  (.A(\vmem[341] ),
    .X(\vmem_after_buf[341] ));
 clkbuf_1 \gen_obs_vmem[342].sdcbuf_gen_vmem  (.A(\vmem[342] ),
    .X(\vmem_after_buf[342] ));
 clkbuf_1 \gen_obs_vmem[343].sdcbuf_gen_vmem  (.A(\vmem[343] ),
    .X(\vmem_after_buf[343] ));
 clkbuf_1 \gen_obs_vmem[344].sdcbuf_gen_vmem  (.A(\vmem[344] ),
    .X(\vmem_after_buf[344] ));
 clkbuf_1 \gen_obs_vmem[345].sdcbuf_gen_vmem  (.A(\vmem[345] ),
    .X(\vmem_after_buf[345] ));
 clkbuf_1 \gen_obs_vmem[346].sdcbuf_gen_vmem  (.A(\vmem[346] ),
    .X(\vmem_after_buf[346] ));
 clkbuf_1 \gen_obs_vmem[347].sdcbuf_gen_vmem  (.A(\vmem[347] ),
    .X(\vmem_after_buf[347] ));
 clkbuf_1 \gen_obs_vmem[348].sdcbuf_gen_vmem  (.A(\vmem[348] ),
    .X(\vmem_after_buf[348] ));
 clkbuf_1 \gen_obs_vmem[349].sdcbuf_gen_vmem  (.A(\vmem[349] ),
    .X(\vmem_after_buf[349] ));
 clkbuf_1 \gen_obs_vmem[34].sdcbuf_gen_vmem  (.A(\vmem[34] ),
    .X(\vmem_after_buf[34] ));
 clkbuf_1 \gen_obs_vmem[350].sdcbuf_gen_vmem  (.A(\vmem[350] ),
    .X(\vmem_after_buf[350] ));
 clkbuf_1 \gen_obs_vmem[351].sdcbuf_gen_vmem  (.A(\vmem[351] ),
    .X(\vmem_after_buf[351] ));
 clkbuf_1 \gen_obs_vmem[352].sdcbuf_gen_vmem  (.A(\vmem[352] ),
    .X(\vmem_after_buf[352] ));
 clkbuf_1 \gen_obs_vmem[353].sdcbuf_gen_vmem  (.A(\vmem[353] ),
    .X(\vmem_after_buf[353] ));
 clkbuf_1 \gen_obs_vmem[354].sdcbuf_gen_vmem  (.A(\vmem[354] ),
    .X(\vmem_after_buf[354] ));
 clkbuf_1 \gen_obs_vmem[355].sdcbuf_gen_vmem  (.A(\vmem[355] ),
    .X(\vmem_after_buf[355] ));
 clkbuf_1 \gen_obs_vmem[356].sdcbuf_gen_vmem  (.A(\vmem[356] ),
    .X(\vmem_after_buf[356] ));
 clkbuf_1 \gen_obs_vmem[357].sdcbuf_gen_vmem  (.A(\vmem[357] ),
    .X(\vmem_after_buf[357] ));
 clkbuf_1 \gen_obs_vmem[358].sdcbuf_gen_vmem  (.A(\vmem[358] ),
    .X(\vmem_after_buf[358] ));
 clkbuf_1 \gen_obs_vmem[359].sdcbuf_gen_vmem  (.A(\vmem[359] ),
    .X(\vmem_after_buf[359] ));
 clkbuf_1 \gen_obs_vmem[35].sdcbuf_gen_vmem  (.A(\vmem[35] ),
    .X(\vmem_after_buf[35] ));
 clkbuf_1 \gen_obs_vmem[360].sdcbuf_gen_vmem  (.A(\vmem[360] ),
    .X(\vmem_after_buf[360] ));
 clkbuf_1 \gen_obs_vmem[361].sdcbuf_gen_vmem  (.A(\vmem[361] ),
    .X(\vmem_after_buf[361] ));
 clkbuf_1 \gen_obs_vmem[362].sdcbuf_gen_vmem  (.A(\vmem[362] ),
    .X(\vmem_after_buf[362] ));
 clkbuf_1 \gen_obs_vmem[363].sdcbuf_gen_vmem  (.A(\vmem[363] ),
    .X(\vmem_after_buf[363] ));
 clkbuf_1 \gen_obs_vmem[364].sdcbuf_gen_vmem  (.A(\vmem[364] ),
    .X(\vmem_after_buf[364] ));
 clkbuf_1 \gen_obs_vmem[365].sdcbuf_gen_vmem  (.A(\vmem[365] ),
    .X(\vmem_after_buf[365] ));
 clkbuf_1 \gen_obs_vmem[366].sdcbuf_gen_vmem  (.A(\vmem[366] ),
    .X(\vmem_after_buf[366] ));
 clkbuf_1 \gen_obs_vmem[367].sdcbuf_gen_vmem  (.A(\vmem[367] ),
    .X(\vmem_after_buf[367] ));
 clkbuf_1 \gen_obs_vmem[368].sdcbuf_gen_vmem  (.A(\vmem[368] ),
    .X(\vmem_after_buf[368] ));
 clkbuf_1 \gen_obs_vmem[369].sdcbuf_gen_vmem  (.A(\vmem[369] ),
    .X(\vmem_after_buf[369] ));
 clkbuf_1 \gen_obs_vmem[36].sdcbuf_gen_vmem  (.A(\vmem[36] ),
    .X(\vmem_after_buf[36] ));
 clkbuf_1 \gen_obs_vmem[370].sdcbuf_gen_vmem  (.A(\vmem[370] ),
    .X(\vmem_after_buf[370] ));
 clkbuf_1 \gen_obs_vmem[371].sdcbuf_gen_vmem  (.A(\vmem[371] ),
    .X(\vmem_after_buf[371] ));
 clkbuf_1 \gen_obs_vmem[372].sdcbuf_gen_vmem  (.A(\vmem[372] ),
    .X(\vmem_after_buf[372] ));
 clkbuf_1 \gen_obs_vmem[373].sdcbuf_gen_vmem  (.A(\vmem[373] ),
    .X(\vmem_after_buf[373] ));
 clkbuf_1 \gen_obs_vmem[374].sdcbuf_gen_vmem  (.A(\vmem[374] ),
    .X(\vmem_after_buf[374] ));
 clkbuf_1 \gen_obs_vmem[375].sdcbuf_gen_vmem  (.A(\vmem[375] ),
    .X(\vmem_after_buf[375] ));
 clkbuf_1 \gen_obs_vmem[376].sdcbuf_gen_vmem  (.A(\vmem[376] ),
    .X(\vmem_after_buf[376] ));
 clkbuf_1 \gen_obs_vmem[377].sdcbuf_gen_vmem  (.A(\vmem[377] ),
    .X(\vmem_after_buf[377] ));
 clkbuf_1 \gen_obs_vmem[378].sdcbuf_gen_vmem  (.A(\vmem[378] ),
    .X(\vmem_after_buf[378] ));
 clkbuf_1 \gen_obs_vmem[379].sdcbuf_gen_vmem  (.A(\vmem[379] ),
    .X(\vmem_after_buf[379] ));
 clkbuf_1 \gen_obs_vmem[37].sdcbuf_gen_vmem  (.A(\vmem[37] ),
    .X(\vmem_after_buf[37] ));
 clkbuf_1 \gen_obs_vmem[380].sdcbuf_gen_vmem  (.A(\vmem[380] ),
    .X(\vmem_after_buf[380] ));
 clkbuf_1 \gen_obs_vmem[381].sdcbuf_gen_vmem  (.A(\vmem[381] ),
    .X(\vmem_after_buf[381] ));
 clkbuf_1 \gen_obs_vmem[382].sdcbuf_gen_vmem  (.A(\vmem[382] ),
    .X(\vmem_after_buf[382] ));
 clkbuf_1 \gen_obs_vmem[383].sdcbuf_gen_vmem  (.A(\vmem[383] ),
    .X(\vmem_after_buf[383] ));
 clkbuf_1 \gen_obs_vmem[384].sdcbuf_gen_vmem  (.A(\vmem[384] ),
    .X(\vmem_after_buf[384] ));
 clkbuf_1 \gen_obs_vmem[385].sdcbuf_gen_vmem  (.A(\vmem[385] ),
    .X(\vmem_after_buf[385] ));
 clkbuf_1 \gen_obs_vmem[386].sdcbuf_gen_vmem  (.A(\vmem[386] ),
    .X(\vmem_after_buf[386] ));
 clkbuf_1 \gen_obs_vmem[387].sdcbuf_gen_vmem  (.A(\vmem[387] ),
    .X(\vmem_after_buf[387] ));
 clkbuf_1 \gen_obs_vmem[388].sdcbuf_gen_vmem  (.A(\vmem[388] ),
    .X(\vmem_after_buf[388] ));
 clkbuf_1 \gen_obs_vmem[389].sdcbuf_gen_vmem  (.A(\vmem[389] ),
    .X(\vmem_after_buf[389] ));
 clkbuf_1 \gen_obs_vmem[38].sdcbuf_gen_vmem  (.A(\vmem[38] ),
    .X(\vmem_after_buf[38] ));
 clkbuf_1 \gen_obs_vmem[390].sdcbuf_gen_vmem  (.A(\vmem[390] ),
    .X(\vmem_after_buf[390] ));
 clkbuf_1 \gen_obs_vmem[391].sdcbuf_gen_vmem  (.A(\vmem[391] ),
    .X(\vmem_after_buf[391] ));
 clkbuf_1 \gen_obs_vmem[392].sdcbuf_gen_vmem  (.A(\vmem[392] ),
    .X(\vmem_after_buf[392] ));
 clkbuf_1 \gen_obs_vmem[393].sdcbuf_gen_vmem  (.A(\vmem[393] ),
    .X(\vmem_after_buf[393] ));
 clkbuf_1 \gen_obs_vmem[394].sdcbuf_gen_vmem  (.A(\vmem[394] ),
    .X(\vmem_after_buf[394] ));
 clkbuf_1 \gen_obs_vmem[395].sdcbuf_gen_vmem  (.A(\vmem[395] ),
    .X(\vmem_after_buf[395] ));
 clkbuf_1 \gen_obs_vmem[396].sdcbuf_gen_vmem  (.A(\vmem[396] ),
    .X(\vmem_after_buf[396] ));
 clkbuf_1 \gen_obs_vmem[397].sdcbuf_gen_vmem  (.A(\vmem[397] ),
    .X(\vmem_after_buf[397] ));
 clkbuf_1 \gen_obs_vmem[398].sdcbuf_gen_vmem  (.A(\vmem[398] ),
    .X(\vmem_after_buf[398] ));
 clkbuf_1 \gen_obs_vmem[399].sdcbuf_gen_vmem  (.A(\vmem[399] ),
    .X(\vmem_after_buf[399] ));
 clkbuf_1 \gen_obs_vmem[39].sdcbuf_gen_vmem  (.A(\vmem[39] ),
    .X(\vmem_after_buf[39] ));
 clkbuf_1 \gen_obs_vmem[3].sdcbuf_gen_vmem  (.A(\vmem[3] ),
    .X(\vmem_after_buf[3] ));
 clkbuf_1 \gen_obs_vmem[400].sdcbuf_gen_vmem  (.A(\vmem[400] ),
    .X(\vmem_after_buf[400] ));
 clkbuf_1 \gen_obs_vmem[401].sdcbuf_gen_vmem  (.A(\vmem[401] ),
    .X(\vmem_after_buf[401] ));
 clkbuf_1 \gen_obs_vmem[402].sdcbuf_gen_vmem  (.A(\vmem[402] ),
    .X(\vmem_after_buf[402] ));
 clkbuf_1 \gen_obs_vmem[403].sdcbuf_gen_vmem  (.A(\vmem[403] ),
    .X(\vmem_after_buf[403] ));
 clkbuf_1 \gen_obs_vmem[404].sdcbuf_gen_vmem  (.A(\vmem[404] ),
    .X(\vmem_after_buf[404] ));
 clkbuf_1 \gen_obs_vmem[405].sdcbuf_gen_vmem  (.A(\vmem[405] ),
    .X(\vmem_after_buf[405] ));
 clkbuf_1 \gen_obs_vmem[406].sdcbuf_gen_vmem  (.A(\vmem[406] ),
    .X(\vmem_after_buf[406] ));
 clkbuf_1 \gen_obs_vmem[407].sdcbuf_gen_vmem  (.A(\vmem[407] ),
    .X(\vmem_after_buf[407] ));
 clkbuf_1 \gen_obs_vmem[408].sdcbuf_gen_vmem  (.A(\vmem[408] ),
    .X(\vmem_after_buf[408] ));
 clkbuf_1 \gen_obs_vmem[409].sdcbuf_gen_vmem  (.A(\vmem[409] ),
    .X(\vmem_after_buf[409] ));
 clkbuf_1 \gen_obs_vmem[40].sdcbuf_gen_vmem  (.A(\vmem[40] ),
    .X(\vmem_after_buf[40] ));
 clkbuf_1 \gen_obs_vmem[410].sdcbuf_gen_vmem  (.A(\vmem[410] ),
    .X(\vmem_after_buf[410] ));
 clkbuf_1 \gen_obs_vmem[411].sdcbuf_gen_vmem  (.A(\vmem[411] ),
    .X(\vmem_after_buf[411] ));
 clkbuf_1 \gen_obs_vmem[412].sdcbuf_gen_vmem  (.A(\vmem[412] ),
    .X(\vmem_after_buf[412] ));
 clkbuf_1 \gen_obs_vmem[413].sdcbuf_gen_vmem  (.A(\vmem[413] ),
    .X(\vmem_after_buf[413] ));
 clkbuf_1 \gen_obs_vmem[414].sdcbuf_gen_vmem  (.A(\vmem[414] ),
    .X(\vmem_after_buf[414] ));
 clkbuf_1 \gen_obs_vmem[415].sdcbuf_gen_vmem  (.A(\vmem[415] ),
    .X(\vmem_after_buf[415] ));
 clkbuf_1 \gen_obs_vmem[416].sdcbuf_gen_vmem  (.A(\vmem[416] ),
    .X(\vmem_after_buf[416] ));
 clkbuf_1 \gen_obs_vmem[417].sdcbuf_gen_vmem  (.A(\vmem[417] ),
    .X(\vmem_after_buf[417] ));
 clkbuf_1 \gen_obs_vmem[418].sdcbuf_gen_vmem  (.A(\vmem[418] ),
    .X(\vmem_after_buf[418] ));
 clkbuf_1 \gen_obs_vmem[419].sdcbuf_gen_vmem  (.A(\vmem[419] ),
    .X(\vmem_after_buf[419] ));
 clkbuf_1 \gen_obs_vmem[41].sdcbuf_gen_vmem  (.A(\vmem[41] ),
    .X(\vmem_after_buf[41] ));
 clkbuf_1 \gen_obs_vmem[420].sdcbuf_gen_vmem  (.A(\vmem[420] ),
    .X(\vmem_after_buf[420] ));
 clkbuf_1 \gen_obs_vmem[421].sdcbuf_gen_vmem  (.A(\vmem[421] ),
    .X(\vmem_after_buf[421] ));
 clkbuf_1 \gen_obs_vmem[422].sdcbuf_gen_vmem  (.A(\vmem[422] ),
    .X(\vmem_after_buf[422] ));
 clkbuf_1 \gen_obs_vmem[423].sdcbuf_gen_vmem  (.A(\vmem[423] ),
    .X(\vmem_after_buf[423] ));
 clkbuf_1 \gen_obs_vmem[424].sdcbuf_gen_vmem  (.A(\vmem[424] ),
    .X(\vmem_after_buf[424] ));
 clkbuf_1 \gen_obs_vmem[425].sdcbuf_gen_vmem  (.A(\vmem[425] ),
    .X(\vmem_after_buf[425] ));
 clkbuf_1 \gen_obs_vmem[426].sdcbuf_gen_vmem  (.A(\vmem[426] ),
    .X(\vmem_after_buf[426] ));
 clkbuf_1 \gen_obs_vmem[427].sdcbuf_gen_vmem  (.A(\vmem[427] ),
    .X(\vmem_after_buf[427] ));
 clkbuf_1 \gen_obs_vmem[428].sdcbuf_gen_vmem  (.A(\vmem[428] ),
    .X(\vmem_after_buf[428] ));
 clkbuf_1 \gen_obs_vmem[429].sdcbuf_gen_vmem  (.A(\vmem[429] ),
    .X(\vmem_after_buf[429] ));
 clkbuf_1 \gen_obs_vmem[42].sdcbuf_gen_vmem  (.A(\vmem[42] ),
    .X(\vmem_after_buf[42] ));
 clkbuf_1 \gen_obs_vmem[430].sdcbuf_gen_vmem  (.A(\vmem[430] ),
    .X(\vmem_after_buf[430] ));
 clkbuf_1 \gen_obs_vmem[431].sdcbuf_gen_vmem  (.A(\vmem[431] ),
    .X(\vmem_after_buf[431] ));
 clkbuf_1 \gen_obs_vmem[432].sdcbuf_gen_vmem  (.A(\vmem[432] ),
    .X(\vmem_after_buf[432] ));
 clkbuf_1 \gen_obs_vmem[433].sdcbuf_gen_vmem  (.A(\vmem[433] ),
    .X(\vmem_after_buf[433] ));
 clkbuf_1 \gen_obs_vmem[434].sdcbuf_gen_vmem  (.A(\vmem[434] ),
    .X(\vmem_after_buf[434] ));
 clkbuf_1 \gen_obs_vmem[435].sdcbuf_gen_vmem  (.A(\vmem[435] ),
    .X(\vmem_after_buf[435] ));
 clkbuf_1 \gen_obs_vmem[436].sdcbuf_gen_vmem  (.A(\vmem[436] ),
    .X(\vmem_after_buf[436] ));
 clkbuf_1 \gen_obs_vmem[437].sdcbuf_gen_vmem  (.A(\vmem[437] ),
    .X(\vmem_after_buf[437] ));
 clkbuf_1 \gen_obs_vmem[438].sdcbuf_gen_vmem  (.A(\vmem[438] ),
    .X(\vmem_after_buf[438] ));
 clkbuf_1 \gen_obs_vmem[439].sdcbuf_gen_vmem  (.A(\vmem[439] ),
    .X(\vmem_after_buf[439] ));
 clkbuf_1 \gen_obs_vmem[43].sdcbuf_gen_vmem  (.A(\vmem[43] ),
    .X(\vmem_after_buf[43] ));
 clkbuf_1 \gen_obs_vmem[440].sdcbuf_gen_vmem  (.A(\vmem[440] ),
    .X(\vmem_after_buf[440] ));
 clkbuf_1 \gen_obs_vmem[441].sdcbuf_gen_vmem  (.A(\vmem[441] ),
    .X(\vmem_after_buf[441] ));
 clkbuf_1 \gen_obs_vmem[442].sdcbuf_gen_vmem  (.A(\vmem[442] ),
    .X(\vmem_after_buf[442] ));
 clkbuf_1 \gen_obs_vmem[443].sdcbuf_gen_vmem  (.A(\vmem[443] ),
    .X(\vmem_after_buf[443] ));
 clkbuf_1 \gen_obs_vmem[444].sdcbuf_gen_vmem  (.A(\vmem[444] ),
    .X(\vmem_after_buf[444] ));
 clkbuf_1 \gen_obs_vmem[445].sdcbuf_gen_vmem  (.A(\vmem[445] ),
    .X(\vmem_after_buf[445] ));
 clkbuf_1 \gen_obs_vmem[446].sdcbuf_gen_vmem  (.A(\vmem[446] ),
    .X(\vmem_after_buf[446] ));
 clkbuf_1 \gen_obs_vmem[447].sdcbuf_gen_vmem  (.A(\vmem[447] ),
    .X(\vmem_after_buf[447] ));
 clkbuf_1 \gen_obs_vmem[448].sdcbuf_gen_vmem  (.A(\vmem[448] ),
    .X(\vmem_after_buf[448] ));
 clkbuf_1 \gen_obs_vmem[449].sdcbuf_gen_vmem  (.A(\vmem[449] ),
    .X(\vmem_after_buf[449] ));
 clkbuf_1 \gen_obs_vmem[44].sdcbuf_gen_vmem  (.A(\vmem[44] ),
    .X(\vmem_after_buf[44] ));
 clkbuf_1 \gen_obs_vmem[450].sdcbuf_gen_vmem  (.A(\vmem[450] ),
    .X(\vmem_after_buf[450] ));
 clkbuf_1 \gen_obs_vmem[451].sdcbuf_gen_vmem  (.A(\vmem[451] ),
    .X(\vmem_after_buf[451] ));
 clkbuf_1 \gen_obs_vmem[452].sdcbuf_gen_vmem  (.A(\vmem[452] ),
    .X(\vmem_after_buf[452] ));
 clkbuf_1 \gen_obs_vmem[453].sdcbuf_gen_vmem  (.A(\vmem[453] ),
    .X(\vmem_after_buf[453] ));
 clkbuf_1 \gen_obs_vmem[454].sdcbuf_gen_vmem  (.A(\vmem[454] ),
    .X(\vmem_after_buf[454] ));
 clkbuf_1 \gen_obs_vmem[455].sdcbuf_gen_vmem  (.A(\vmem[455] ),
    .X(\vmem_after_buf[455] ));
 clkbuf_1 \gen_obs_vmem[456].sdcbuf_gen_vmem  (.A(\vmem[456] ),
    .X(\vmem_after_buf[456] ));
 clkbuf_1 \gen_obs_vmem[457].sdcbuf_gen_vmem  (.A(\vmem[457] ),
    .X(\vmem_after_buf[457] ));
 clkbuf_1 \gen_obs_vmem[458].sdcbuf_gen_vmem  (.A(\vmem[458] ),
    .X(\vmem_after_buf[458] ));
 clkbuf_1 \gen_obs_vmem[459].sdcbuf_gen_vmem  (.A(\vmem[459] ),
    .X(\vmem_after_buf[459] ));
 clkbuf_1 \gen_obs_vmem[45].sdcbuf_gen_vmem  (.A(\vmem[45] ),
    .X(\vmem_after_buf[45] ));
 clkbuf_1 \gen_obs_vmem[460].sdcbuf_gen_vmem  (.A(\vmem[460] ),
    .X(\vmem_after_buf[460] ));
 clkbuf_1 \gen_obs_vmem[461].sdcbuf_gen_vmem  (.A(\vmem[461] ),
    .X(\vmem_after_buf[461] ));
 clkbuf_1 \gen_obs_vmem[462].sdcbuf_gen_vmem  (.A(\vmem[462] ),
    .X(\vmem_after_buf[462] ));
 clkbuf_1 \gen_obs_vmem[463].sdcbuf_gen_vmem  (.A(\vmem[463] ),
    .X(\vmem_after_buf[463] ));
 clkbuf_1 \gen_obs_vmem[464].sdcbuf_gen_vmem  (.A(\vmem[464] ),
    .X(\vmem_after_buf[464] ));
 clkbuf_1 \gen_obs_vmem[465].sdcbuf_gen_vmem  (.A(\vmem[465] ),
    .X(\vmem_after_buf[465] ));
 clkbuf_1 \gen_obs_vmem[466].sdcbuf_gen_vmem  (.A(\vmem[466] ),
    .X(\vmem_after_buf[466] ));
 clkbuf_1 \gen_obs_vmem[467].sdcbuf_gen_vmem  (.A(\vmem[467] ),
    .X(\vmem_after_buf[467] ));
 clkbuf_1 \gen_obs_vmem[468].sdcbuf_gen_vmem  (.A(\vmem[468] ),
    .X(\vmem_after_buf[468] ));
 clkbuf_1 \gen_obs_vmem[469].sdcbuf_gen_vmem  (.A(\vmem[469] ),
    .X(\vmem_after_buf[469] ));
 clkbuf_1 \gen_obs_vmem[46].sdcbuf_gen_vmem  (.A(\vmem[46] ),
    .X(\vmem_after_buf[46] ));
 clkbuf_1 \gen_obs_vmem[470].sdcbuf_gen_vmem  (.A(\vmem[470] ),
    .X(\vmem_after_buf[470] ));
 clkbuf_1 \gen_obs_vmem[471].sdcbuf_gen_vmem  (.A(\vmem[471] ),
    .X(\vmem_after_buf[471] ));
 clkbuf_1 \gen_obs_vmem[472].sdcbuf_gen_vmem  (.A(\vmem[472] ),
    .X(\vmem_after_buf[472] ));
 clkbuf_1 \gen_obs_vmem[473].sdcbuf_gen_vmem  (.A(\vmem[473] ),
    .X(\vmem_after_buf[473] ));
 clkbuf_1 \gen_obs_vmem[474].sdcbuf_gen_vmem  (.A(\vmem[474] ),
    .X(\vmem_after_buf[474] ));
 clkbuf_1 \gen_obs_vmem[475].sdcbuf_gen_vmem  (.A(\vmem[475] ),
    .X(\vmem_after_buf[475] ));
 clkbuf_1 \gen_obs_vmem[476].sdcbuf_gen_vmem  (.A(\vmem[476] ),
    .X(\vmem_after_buf[476] ));
 clkbuf_1 \gen_obs_vmem[477].sdcbuf_gen_vmem  (.A(\vmem[477] ),
    .X(\vmem_after_buf[477] ));
 clkbuf_1 \gen_obs_vmem[478].sdcbuf_gen_vmem  (.A(\vmem[478] ),
    .X(\vmem_after_buf[478] ));
 clkbuf_1 \gen_obs_vmem[479].sdcbuf_gen_vmem  (.A(\vmem[479] ),
    .X(\vmem_after_buf[479] ));
 clkbuf_1 \gen_obs_vmem[47].sdcbuf_gen_vmem  (.A(\vmem[47] ),
    .X(\vmem_after_buf[47] ));
 clkbuf_1 \gen_obs_vmem[480].sdcbuf_gen_vmem  (.A(\vmem[480] ),
    .X(\vmem_after_buf[480] ));
 clkbuf_1 \gen_obs_vmem[481].sdcbuf_gen_vmem  (.A(\vmem[481] ),
    .X(\vmem_after_buf[481] ));
 clkbuf_1 \gen_obs_vmem[482].sdcbuf_gen_vmem  (.A(\vmem[482] ),
    .X(\vmem_after_buf[482] ));
 clkbuf_1 \gen_obs_vmem[483].sdcbuf_gen_vmem  (.A(\vmem[483] ),
    .X(\vmem_after_buf[483] ));
 clkbuf_1 \gen_obs_vmem[484].sdcbuf_gen_vmem  (.A(\vmem[484] ),
    .X(\vmem_after_buf[484] ));
 clkbuf_1 \gen_obs_vmem[485].sdcbuf_gen_vmem  (.A(\vmem[485] ),
    .X(\vmem_after_buf[485] ));
 clkbuf_1 \gen_obs_vmem[486].sdcbuf_gen_vmem  (.A(\vmem[486] ),
    .X(\vmem_after_buf[486] ));
 clkbuf_1 \gen_obs_vmem[487].sdcbuf_gen_vmem  (.A(\vmem[487] ),
    .X(\vmem_after_buf[487] ));
 clkbuf_1 \gen_obs_vmem[488].sdcbuf_gen_vmem  (.A(\vmem[488] ),
    .X(\vmem_after_buf[488] ));
 clkbuf_1 \gen_obs_vmem[489].sdcbuf_gen_vmem  (.A(\vmem[489] ),
    .X(\vmem_after_buf[489] ));
 clkbuf_1 \gen_obs_vmem[48].sdcbuf_gen_vmem  (.A(\vmem[48] ),
    .X(\vmem_after_buf[48] ));
 clkbuf_1 \gen_obs_vmem[490].sdcbuf_gen_vmem  (.A(\vmem[490] ),
    .X(\vmem_after_buf[490] ));
 clkbuf_1 \gen_obs_vmem[491].sdcbuf_gen_vmem  (.A(\vmem[491] ),
    .X(\vmem_after_buf[491] ));
 clkbuf_1 \gen_obs_vmem[492].sdcbuf_gen_vmem  (.A(\vmem[492] ),
    .X(\vmem_after_buf[492] ));
 clkbuf_1 \gen_obs_vmem[493].sdcbuf_gen_vmem  (.A(\vmem[493] ),
    .X(\vmem_after_buf[493] ));
 clkbuf_1 \gen_obs_vmem[494].sdcbuf_gen_vmem  (.A(\vmem[494] ),
    .X(\vmem_after_buf[494] ));
 clkbuf_1 \gen_obs_vmem[495].sdcbuf_gen_vmem  (.A(\vmem[495] ),
    .X(\vmem_after_buf[495] ));
 clkbuf_1 \gen_obs_vmem[496].sdcbuf_gen_vmem  (.A(\vmem[496] ),
    .X(\vmem_after_buf[496] ));
 clkbuf_1 \gen_obs_vmem[497].sdcbuf_gen_vmem  (.A(\vmem[497] ),
    .X(\vmem_after_buf[497] ));
 clkbuf_1 \gen_obs_vmem[498].sdcbuf_gen_vmem  (.A(\vmem[498] ),
    .X(\vmem_after_buf[498] ));
 clkbuf_1 \gen_obs_vmem[499].sdcbuf_gen_vmem  (.A(\vmem[499] ),
    .X(\vmem_after_buf[499] ));
 clkbuf_1 \gen_obs_vmem[49].sdcbuf_gen_vmem  (.A(\vmem[49] ),
    .X(\vmem_after_buf[49] ));
 clkbuf_1 \gen_obs_vmem[4].sdcbuf_gen_vmem  (.A(\vmem[4] ),
    .X(\vmem_after_buf[4] ));
 clkbuf_1 \gen_obs_vmem[500].sdcbuf_gen_vmem  (.A(\vmem[500] ),
    .X(\vmem_after_buf[500] ));
 clkbuf_1 \gen_obs_vmem[501].sdcbuf_gen_vmem  (.A(\vmem[501] ),
    .X(\vmem_after_buf[501] ));
 clkbuf_1 \gen_obs_vmem[502].sdcbuf_gen_vmem  (.A(\vmem[502] ),
    .X(\vmem_after_buf[502] ));
 clkbuf_1 \gen_obs_vmem[503].sdcbuf_gen_vmem  (.A(\vmem[503] ),
    .X(\vmem_after_buf[503] ));
 clkbuf_1 \gen_obs_vmem[504].sdcbuf_gen_vmem  (.A(\vmem[504] ),
    .X(\vmem_after_buf[504] ));
 clkbuf_1 \gen_obs_vmem[505].sdcbuf_gen_vmem  (.A(\vmem[505] ),
    .X(\vmem_after_buf[505] ));
 clkbuf_1 \gen_obs_vmem[506].sdcbuf_gen_vmem  (.A(\vmem[506] ),
    .X(\vmem_after_buf[506] ));
 clkbuf_1 \gen_obs_vmem[507].sdcbuf_gen_vmem  (.A(\vmem[507] ),
    .X(\vmem_after_buf[507] ));
 clkbuf_1 \gen_obs_vmem[508].sdcbuf_gen_vmem  (.A(\vmem[508] ),
    .X(\vmem_after_buf[508] ));
 clkbuf_1 \gen_obs_vmem[509].sdcbuf_gen_vmem  (.A(\vmem[509] ),
    .X(\vmem_after_buf[509] ));
 clkbuf_1 \gen_obs_vmem[50].sdcbuf_gen_vmem  (.A(\vmem[50] ),
    .X(\vmem_after_buf[50] ));
 clkbuf_1 \gen_obs_vmem[510].sdcbuf_gen_vmem  (.A(\vmem[510] ),
    .X(\vmem_after_buf[510] ));
 clkbuf_1 \gen_obs_vmem[511].sdcbuf_gen_vmem  (.A(\vmem[511] ),
    .X(\vmem_after_buf[511] ));
 clkbuf_1 \gen_obs_vmem[51].sdcbuf_gen_vmem  (.A(\vmem[51] ),
    .X(\vmem_after_buf[51] ));
 clkbuf_1 \gen_obs_vmem[52].sdcbuf_gen_vmem  (.A(\vmem[52] ),
    .X(\vmem_after_buf[52] ));
 clkbuf_1 \gen_obs_vmem[53].sdcbuf_gen_vmem  (.A(\vmem[53] ),
    .X(\vmem_after_buf[53] ));
 clkbuf_1 \gen_obs_vmem[54].sdcbuf_gen_vmem  (.A(\vmem[54] ),
    .X(\vmem_after_buf[54] ));
 clkbuf_1 \gen_obs_vmem[55].sdcbuf_gen_vmem  (.A(\vmem[55] ),
    .X(\vmem_after_buf[55] ));
 clkbuf_1 \gen_obs_vmem[56].sdcbuf_gen_vmem  (.A(\vmem[56] ),
    .X(\vmem_after_buf[56] ));
 clkbuf_1 \gen_obs_vmem[57].sdcbuf_gen_vmem  (.A(\vmem[57] ),
    .X(\vmem_after_buf[57] ));
 clkbuf_1 \gen_obs_vmem[58].sdcbuf_gen_vmem  (.A(\vmem[58] ),
    .X(\vmem_after_buf[58] ));
 clkbuf_1 \gen_obs_vmem[59].sdcbuf_gen_vmem  (.A(\vmem[59] ),
    .X(\vmem_after_buf[59] ));
 clkbuf_1 \gen_obs_vmem[5].sdcbuf_gen_vmem  (.A(\vmem[5] ),
    .X(\vmem_after_buf[5] ));
 clkbuf_1 \gen_obs_vmem[60].sdcbuf_gen_vmem  (.A(\vmem[60] ),
    .X(\vmem_after_buf[60] ));
 clkbuf_1 \gen_obs_vmem[61].sdcbuf_gen_vmem  (.A(\vmem[61] ),
    .X(\vmem_after_buf[61] ));
 clkbuf_1 \gen_obs_vmem[62].sdcbuf_gen_vmem  (.A(\vmem[62] ),
    .X(\vmem_after_buf[62] ));
 clkbuf_1 \gen_obs_vmem[63].sdcbuf_gen_vmem  (.A(\vmem[63] ),
    .X(\vmem_after_buf[63] ));
 clkbuf_1 \gen_obs_vmem[64].sdcbuf_gen_vmem  (.A(\vmem[64] ),
    .X(\vmem_after_buf[64] ));
 clkbuf_1 \gen_obs_vmem[65].sdcbuf_gen_vmem  (.A(\vmem[65] ),
    .X(\vmem_after_buf[65] ));
 clkbuf_1 \gen_obs_vmem[66].sdcbuf_gen_vmem  (.A(\vmem[66] ),
    .X(\vmem_after_buf[66] ));
 clkbuf_1 \gen_obs_vmem[67].sdcbuf_gen_vmem  (.A(\vmem[67] ),
    .X(\vmem_after_buf[67] ));
 clkbuf_1 \gen_obs_vmem[68].sdcbuf_gen_vmem  (.A(\vmem[68] ),
    .X(\vmem_after_buf[68] ));
 clkbuf_1 \gen_obs_vmem[69].sdcbuf_gen_vmem  (.A(\vmem[69] ),
    .X(\vmem_after_buf[69] ));
 clkbuf_1 \gen_obs_vmem[6].sdcbuf_gen_vmem  (.A(\vmem[6] ),
    .X(\vmem_after_buf[6] ));
 clkbuf_1 \gen_obs_vmem[70].sdcbuf_gen_vmem  (.A(\vmem[70] ),
    .X(\vmem_after_buf[70] ));
 clkbuf_1 \gen_obs_vmem[71].sdcbuf_gen_vmem  (.A(\vmem[71] ),
    .X(\vmem_after_buf[71] ));
 clkbuf_1 \gen_obs_vmem[72].sdcbuf_gen_vmem  (.A(\vmem[72] ),
    .X(\vmem_after_buf[72] ));
 clkbuf_1 \gen_obs_vmem[73].sdcbuf_gen_vmem  (.A(\vmem[73] ),
    .X(\vmem_after_buf[73] ));
 clkbuf_1 \gen_obs_vmem[74].sdcbuf_gen_vmem  (.A(\vmem[74] ),
    .X(\vmem_after_buf[74] ));
 clkbuf_1 \gen_obs_vmem[75].sdcbuf_gen_vmem  (.A(\vmem[75] ),
    .X(\vmem_after_buf[75] ));
 clkbuf_1 \gen_obs_vmem[76].sdcbuf_gen_vmem  (.A(\vmem[76] ),
    .X(\vmem_after_buf[76] ));
 clkbuf_1 \gen_obs_vmem[77].sdcbuf_gen_vmem  (.A(\vmem[77] ),
    .X(\vmem_after_buf[77] ));
 clkbuf_1 \gen_obs_vmem[78].sdcbuf_gen_vmem  (.A(\vmem[78] ),
    .X(\vmem_after_buf[78] ));
 clkbuf_1 \gen_obs_vmem[79].sdcbuf_gen_vmem  (.A(\vmem[79] ),
    .X(\vmem_after_buf[79] ));
 clkbuf_1 \gen_obs_vmem[7].sdcbuf_gen_vmem  (.A(\vmem[7] ),
    .X(\vmem_after_buf[7] ));
 clkbuf_1 \gen_obs_vmem[80].sdcbuf_gen_vmem  (.A(\vmem[80] ),
    .X(\vmem_after_buf[80] ));
 clkbuf_1 \gen_obs_vmem[81].sdcbuf_gen_vmem  (.A(\vmem[81] ),
    .X(\vmem_after_buf[81] ));
 clkbuf_1 \gen_obs_vmem[82].sdcbuf_gen_vmem  (.A(\vmem[82] ),
    .X(\vmem_after_buf[82] ));
 clkbuf_1 \gen_obs_vmem[83].sdcbuf_gen_vmem  (.A(\vmem[83] ),
    .X(\vmem_after_buf[83] ));
 clkbuf_1 \gen_obs_vmem[84].sdcbuf_gen_vmem  (.A(\vmem[84] ),
    .X(\vmem_after_buf[84] ));
 clkbuf_1 \gen_obs_vmem[85].sdcbuf_gen_vmem  (.A(\vmem[85] ),
    .X(\vmem_after_buf[85] ));
 clkbuf_1 \gen_obs_vmem[86].sdcbuf_gen_vmem  (.A(\vmem[86] ),
    .X(\vmem_after_buf[86] ));
 clkbuf_1 \gen_obs_vmem[87].sdcbuf_gen_vmem  (.A(\vmem[87] ),
    .X(\vmem_after_buf[87] ));
 clkbuf_1 \gen_obs_vmem[88].sdcbuf_gen_vmem  (.A(\vmem[88] ),
    .X(\vmem_after_buf[88] ));
 clkbuf_1 \gen_obs_vmem[89].sdcbuf_gen_vmem  (.A(\vmem[89] ),
    .X(\vmem_after_buf[89] ));
 clkbuf_1 \gen_obs_vmem[8].sdcbuf_gen_vmem  (.A(\vmem[8] ),
    .X(\vmem_after_buf[8] ));
 clkbuf_1 \gen_obs_vmem[90].sdcbuf_gen_vmem  (.A(\vmem[90] ),
    .X(\vmem_after_buf[90] ));
 clkbuf_1 \gen_obs_vmem[91].sdcbuf_gen_vmem  (.A(\vmem[91] ),
    .X(\vmem_after_buf[91] ));
 clkbuf_1 \gen_obs_vmem[92].sdcbuf_gen_vmem  (.A(\vmem[92] ),
    .X(\vmem_after_buf[92] ));
 clkbuf_1 \gen_obs_vmem[93].sdcbuf_gen_vmem  (.A(\vmem[93] ),
    .X(\vmem_after_buf[93] ));
 clkbuf_1 \gen_obs_vmem[94].sdcbuf_gen_vmem  (.A(\vmem[94] ),
    .X(\vmem_after_buf[94] ));
 clkbuf_1 \gen_obs_vmem[95].sdcbuf_gen_vmem  (.A(\vmem[95] ),
    .X(\vmem_after_buf[95] ));
 clkbuf_1 \gen_obs_vmem[96].sdcbuf_gen_vmem  (.A(\vmem[96] ),
    .X(\vmem_after_buf[96] ));
 clkbuf_1 \gen_obs_vmem[97].sdcbuf_gen_vmem  (.A(\vmem[97] ),
    .X(\vmem_after_buf[97] ));
 clkbuf_1 \gen_obs_vmem[98].sdcbuf_gen_vmem  (.A(\vmem[98] ),
    .X(\vmem_after_buf[98] ));
 clkbuf_1 \gen_obs_vmem[99].sdcbuf_gen_vmem  (.A(\vmem[99] ),
    .X(\vmem_after_buf[99] ));
 clkbuf_1 \gen_obs_vmem[9].sdcbuf_gen_vmem  (.A(\vmem[9] ),
    .X(\vmem_after_buf[9] ));
 clkbuf_1 sdcbuf_ff_erase (.A(ff_erase),
    .X(ff_erase_after_buf));
 clkbuf_1 sdcbuf_ff_prog (.A(ff_prog),
    .X(ff_prog_after_buf));
 clkbuf_1 sdcbuf_s1_rst (.A(\digitop_pav2.invent_inst.s1_r_o ),
    .X(s1_rst_after_buf));
 clkbuf_1 sdcbuf_s1_set (.A(\digitop_pav2.invent_inst.s1_s_o ),
    .X(s1_set_after_buf));
 clkbuf_1 sdcbuf_s2_rst (.A(\digitop_pav2.invent_inst.s2_r_o ),
    .X(s2_rst_after_buf));
 clkbuf_1 sdcbuf_s2_set (.A(\digitop_pav2.invent_inst.s2_s_o ),
    .X(s2_set_after_buf));
 clkbuf_1 sdcbuf_s3_rst (.A(\digitop_pav2.invent_inst.s3_r_o ),
    .X(s3_rst_after_buf));
 clkbuf_1 sdcbuf_s3_set (.A(\digitop_pav2.invent_inst.s3_s_o ),
    .X(s3_set_after_buf));
 clkbuf_1 sdcbuf_sl_rst (.A(\digitop_pav2.invent_inst.sl_r_o ),
    .X(sl_rst_after_buf));
 clkbuf_1 sdcbuf_sl_set (.A(\digitop_pav2.invent_inst.sl_s_o ),
    .X(sl_set_after_buf));
 dlygate4sd3_1 \stadly_mpw03_erase_rise_0.stdinst_dlygate4sd3_1  (.A(ff_erase_rise),
    .X(\stadly_mpw03_erase_rise_0.Y ));
 dlygate4sd3_1 \stadly_mpw03_erase_rise_1.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_erase_rise_0.Y ),
    .X(\stadly_mpw03_erase_rise_1.Y ));
 dlygate4sd3_1 \stadly_mpw03_erase_rise_2.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_erase_rise_1.Y ),
    .X(\stadly_mpw03_erase_rise_2.Y ));
 dlygate4sd3_1 \stadly_mpw03_erase_rise_3.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_erase_rise_2.Y ),
    .X(\stadly_mpw03_erase_rise_3.Y ));
 dlygate4sd3_1 \stadly_mpw03_erase_rise_4.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_erase_rise_3.Y ),
    .X(\stadly_mpw03_erase_rise_4.Y ));
 dlygate4sd3_1 \stadly_mpw03_erase_rise_5.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_erase_rise_4.Y ),
    .X(\stadly_mpw03_erase_rise_5.Y ));
 dlygate4sd3_1 \stadly_mpw03_erase_rise_6.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_erase_rise_5.Y ),
    .X(\stadly_mpw03_erase_rise_6.Y ));
 dlygate4sd3_1 \stadly_mpw03_erase_rise_7.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_erase_rise_6.Y ),
    .X(\stadly_mpw03_erase_rise_7.Y ));
 dlygate4sd3_1 \stadly_mpw03_erase_rise_8.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_erase_rise_7.Y ),
    .X(\stadly_mpw03_erase_rise_8.Y ));
 clkbuf_2 \stadly_mpw03_erase_rise_9.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_erase_rise_8.Y ),
    .X(\stadly_mpw03_erase_rise_9.Y ));
 dlygate4sd3_1 \stadly_mpw03_prog_rise_0.stdinst_dlygate4sd3_1  (.A(ff_prog_rise),
    .X(\stadly_mpw03_prog_rise_0.Y ));
 dlygate4sd3_1 \stadly_mpw03_prog_rise_1.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_prog_rise_0.Y ),
    .X(\stadly_mpw03_prog_rise_1.Y ));
 dlygate4sd3_1 \stadly_mpw03_prog_rise_2.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_prog_rise_1.Y ),
    .X(\stadly_mpw03_prog_rise_2.Y ));
 dlygate4sd3_1 \stadly_mpw03_prog_rise_3.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_prog_rise_2.Y ),
    .X(\stadly_mpw03_prog_rise_3.Y ));
 dlygate4sd3_1 \stadly_mpw03_prog_rise_4.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_prog_rise_3.Y ),
    .X(\stadly_mpw03_prog_rise_4.Y ));
 dlygate4sd3_1 \stadly_mpw03_prog_rise_5.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_prog_rise_4.Y ),
    .X(\stadly_mpw03_prog_rise_5.Y ));
 dlygate4sd3_1 \stadly_mpw03_prog_rise_6.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_prog_rise_5.Y ),
    .X(\stadly_mpw03_prog_rise_6.Y ));
 dlygate4sd3_1 \stadly_mpw03_prog_rise_7.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_prog_rise_6.Y ),
    .X(\stadly_mpw03_prog_rise_7.Y ));
 dlygate4sd3_1 \stadly_mpw03_prog_rise_8.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_prog_rise_7.Y ),
    .X(\stadly_mpw03_prog_rise_8.Y ));
 clkbuf_2 \stadly_mpw03_prog_rise_9.stdinst_dlygate4sd3_1  (.A(\stadly_mpw03_prog_rise_8.Y ),
    .X(\stadly_mpw03_prog_rise_9.Y ));
 decap_3 PHY_EDGE_ROW_0_Right_0 ();
 decap_3 PHY_EDGE_ROW_1_Right_1 ();
 decap_3 PHY_EDGE_ROW_2_Right_2 ();
 decap_3 PHY_EDGE_ROW_3_Right_3 ();
 decap_3 PHY_EDGE_ROW_4_Right_4 ();
 decap_3 PHY_EDGE_ROW_5_Right_5 ();
 decap_3 PHY_EDGE_ROW_6_Right_6 ();
 decap_3 PHY_EDGE_ROW_7_Right_7 ();
 decap_3 PHY_EDGE_ROW_8_Right_8 ();
 decap_3 PHY_EDGE_ROW_9_Right_9 ();
 decap_3 PHY_EDGE_ROW_10_Right_10 ();
 decap_3 PHY_EDGE_ROW_11_Right_11 ();
 decap_3 PHY_EDGE_ROW_12_Right_12 ();
 decap_3 PHY_EDGE_ROW_13_Right_13 ();
 decap_3 PHY_EDGE_ROW_14_Right_14 ();
 decap_3 PHY_EDGE_ROW_15_Right_15 ();
 decap_3 PHY_EDGE_ROW_16_Right_16 ();
 decap_3 PHY_EDGE_ROW_17_Right_17 ();
 decap_3 PHY_EDGE_ROW_18_Right_18 ();
 decap_3 PHY_EDGE_ROW_19_Right_19 ();
 decap_3 PHY_EDGE_ROW_20_Right_20 ();
 decap_3 PHY_EDGE_ROW_21_Right_21 ();
 decap_3 PHY_EDGE_ROW_22_Right_22 ();
 decap_3 PHY_EDGE_ROW_23_Right_23 ();
 decap_3 PHY_EDGE_ROW_24_Right_24 ();
 decap_3 PHY_EDGE_ROW_25_Right_25 ();
 decap_3 PHY_EDGE_ROW_26_Right_26 ();
 decap_3 PHY_EDGE_ROW_27_Right_27 ();
 decap_3 PHY_EDGE_ROW_28_Right_28 ();
 decap_3 PHY_EDGE_ROW_29_Right_29 ();
 decap_3 PHY_EDGE_ROW_30_Right_30 ();
 decap_3 PHY_EDGE_ROW_31_Right_31 ();
 decap_3 PHY_EDGE_ROW_32_Right_32 ();
 decap_3 PHY_EDGE_ROW_33_Right_33 ();
 decap_3 PHY_EDGE_ROW_34_Right_34 ();
 decap_3 PHY_EDGE_ROW_35_Right_35 ();
 decap_3 PHY_EDGE_ROW_36_Right_36 ();
 decap_3 PHY_EDGE_ROW_37_Right_37 ();
 decap_3 PHY_EDGE_ROW_38_Right_38 ();
 decap_3 PHY_EDGE_ROW_39_Right_39 ();
 decap_3 PHY_EDGE_ROW_40_Right_40 ();
 decap_3 PHY_EDGE_ROW_41_Right_41 ();
 decap_3 PHY_EDGE_ROW_42_Right_42 ();
 decap_3 PHY_EDGE_ROW_43_Right_43 ();
 decap_3 PHY_EDGE_ROW_44_Right_44 ();
 decap_3 PHY_EDGE_ROW_45_Right_45 ();
 decap_3 PHY_EDGE_ROW_46_Right_46 ();
 decap_3 PHY_EDGE_ROW_47_Right_47 ();
 decap_3 PHY_EDGE_ROW_48_Right_48 ();
 decap_3 PHY_EDGE_ROW_49_Right_49 ();
 decap_3 PHY_EDGE_ROW_50_Right_50 ();
 decap_3 PHY_EDGE_ROW_51_Right_51 ();
 decap_3 PHY_EDGE_ROW_52_Right_52 ();
 decap_3 PHY_EDGE_ROW_53_Right_53 ();
 decap_3 PHY_EDGE_ROW_54_Right_54 ();
 decap_3 PHY_EDGE_ROW_55_Right_55 ();
 decap_3 PHY_EDGE_ROW_56_Right_56 ();
 decap_3 PHY_EDGE_ROW_57_Right_57 ();
 decap_3 PHY_EDGE_ROW_58_Right_58 ();
 decap_3 PHY_EDGE_ROW_59_Right_59 ();
 decap_3 PHY_EDGE_ROW_60_Right_60 ();
 decap_3 PHY_EDGE_ROW_61_Right_61 ();
 decap_3 PHY_EDGE_ROW_62_Right_62 ();
 decap_3 PHY_EDGE_ROW_63_Right_63 ();
 decap_3 PHY_EDGE_ROW_64_Right_64 ();
 decap_3 PHY_EDGE_ROW_65_Right_65 ();
 decap_3 PHY_EDGE_ROW_66_Right_66 ();
 decap_3 PHY_EDGE_ROW_67_Right_67 ();
 decap_3 PHY_EDGE_ROW_68_Right_68 ();
 decap_3 PHY_EDGE_ROW_69_Right_69 ();
 decap_3 PHY_EDGE_ROW_70_Right_70 ();
 decap_3 PHY_EDGE_ROW_71_Right_71 ();
 decap_3 PHY_EDGE_ROW_72_Right_72 ();
 decap_3 PHY_EDGE_ROW_73_Right_73 ();
 decap_3 PHY_EDGE_ROW_74_Right_74 ();
 decap_3 PHY_EDGE_ROW_75_Right_75 ();
 decap_3 PHY_EDGE_ROW_76_Right_76 ();
 decap_3 PHY_EDGE_ROW_77_Right_77 ();
 decap_3 PHY_EDGE_ROW_78_Right_78 ();
 decap_3 PHY_EDGE_ROW_79_Right_79 ();
 decap_3 PHY_EDGE_ROW_80_Right_80 ();
 decap_3 PHY_EDGE_ROW_81_Right_81 ();
 decap_3 PHY_EDGE_ROW_82_Right_82 ();
 decap_3 PHY_EDGE_ROW_83_Right_83 ();
 decap_3 PHY_EDGE_ROW_84_Right_84 ();
 decap_3 PHY_EDGE_ROW_85_Right_85 ();
 decap_3 PHY_EDGE_ROW_86_Right_86 ();
 decap_3 PHY_EDGE_ROW_87_Right_87 ();
 decap_3 PHY_EDGE_ROW_88_Right_88 ();
 decap_3 PHY_EDGE_ROW_89_Right_89 ();
 decap_3 PHY_EDGE_ROW_90_Right_90 ();
 decap_3 PHY_EDGE_ROW_91_Right_91 ();
 decap_3 PHY_EDGE_ROW_92_Right_92 ();
 decap_3 PHY_EDGE_ROW_93_Right_93 ();
 decap_3 PHY_EDGE_ROW_94_Right_94 ();
 decap_3 PHY_EDGE_ROW_95_Right_95 ();
 decap_3 PHY_EDGE_ROW_96_Right_96 ();
 decap_3 PHY_EDGE_ROW_97_Right_97 ();
 decap_3 PHY_EDGE_ROW_98_Right_98 ();
 decap_3 PHY_EDGE_ROW_99_Right_99 ();
 decap_3 PHY_EDGE_ROW_100_Right_100 ();
 decap_3 PHY_EDGE_ROW_101_Right_101 ();
 decap_3 PHY_EDGE_ROW_102_Right_102 ();
 decap_3 PHY_EDGE_ROW_103_Right_103 ();
 decap_3 PHY_EDGE_ROW_104_Right_104 ();
 decap_3 PHY_EDGE_ROW_105_Right_105 ();
 decap_3 PHY_EDGE_ROW_106_Right_106 ();
 decap_3 PHY_EDGE_ROW_107_Right_107 ();
 decap_3 PHY_EDGE_ROW_108_Right_108 ();
 decap_3 PHY_EDGE_ROW_109_Right_109 ();
 decap_3 PHY_EDGE_ROW_110_Right_110 ();
 decap_3 PHY_EDGE_ROW_111_Right_111 ();
 decap_3 PHY_EDGE_ROW_112_Right_112 ();
 decap_3 PHY_EDGE_ROW_113_Right_113 ();
 decap_3 PHY_EDGE_ROW_114_Right_114 ();
 decap_3 PHY_EDGE_ROW_115_Right_115 ();
 decap_3 PHY_EDGE_ROW_116_Right_116 ();
 decap_3 PHY_EDGE_ROW_117_Right_117 ();
 decap_3 PHY_EDGE_ROW_118_Right_118 ();
 decap_3 PHY_EDGE_ROW_119_Right_119 ();
 decap_3 PHY_EDGE_ROW_120_Right_120 ();
 decap_3 PHY_EDGE_ROW_121_Right_121 ();
 decap_3 PHY_EDGE_ROW_122_Right_122 ();
 decap_3 PHY_EDGE_ROW_123_Right_123 ();
 decap_3 PHY_EDGE_ROW_124_Right_124 ();
 decap_3 PHY_EDGE_ROW_125_Right_125 ();
 decap_3 PHY_EDGE_ROW_126_Right_126 ();
 decap_3 PHY_EDGE_ROW_127_Right_127 ();
 decap_3 PHY_EDGE_ROW_128_Right_128 ();
 decap_3 PHY_EDGE_ROW_129_Right_129 ();
 decap_3 PHY_EDGE_ROW_130_Right_130 ();
 decap_3 PHY_EDGE_ROW_131_Right_131 ();
 decap_3 PHY_EDGE_ROW_132_Right_132 ();
 decap_3 PHY_EDGE_ROW_133_Right_133 ();
 decap_3 PHY_EDGE_ROW_134_Right_134 ();
 decap_3 PHY_EDGE_ROW_135_Right_135 ();
 decap_3 PHY_EDGE_ROW_136_Right_136 ();
 decap_3 PHY_EDGE_ROW_137_Right_137 ();
 decap_3 PHY_EDGE_ROW_138_Right_138 ();
 decap_3 PHY_EDGE_ROW_139_Right_139 ();
 decap_3 PHY_EDGE_ROW_140_Right_140 ();
 decap_3 PHY_EDGE_ROW_141_Right_141 ();
 decap_3 PHY_EDGE_ROW_142_Right_142 ();
 decap_3 PHY_EDGE_ROW_143_Right_143 ();
 decap_3 PHY_EDGE_ROW_144_Right_144 ();
 decap_3 PHY_EDGE_ROW_145_Right_145 ();
 decap_3 PHY_EDGE_ROW_146_Right_146 ();
 decap_3 PHY_EDGE_ROW_147_Right_147 ();
 decap_3 PHY_EDGE_ROW_148_Right_148 ();
 decap_3 PHY_EDGE_ROW_149_Right_149 ();
 decap_3 PHY_EDGE_ROW_150_Right_150 ();
 decap_3 PHY_EDGE_ROW_151_Right_151 ();
 decap_3 PHY_EDGE_ROW_152_Right_152 ();
 decap_3 PHY_EDGE_ROW_153_Right_153 ();
 decap_3 PHY_EDGE_ROW_154_Right_154 ();
 decap_3 PHY_EDGE_ROW_155_Right_155 ();
 decap_3 PHY_EDGE_ROW_156_Right_156 ();
 decap_3 PHY_EDGE_ROW_157_Right_157 ();
 decap_3 PHY_EDGE_ROW_158_Right_158 ();
 decap_3 PHY_EDGE_ROW_159_Right_159 ();
 decap_3 PHY_EDGE_ROW_160_Right_160 ();
 decap_3 PHY_EDGE_ROW_161_Right_161 ();
 decap_3 PHY_EDGE_ROW_162_Right_162 ();
 decap_3 PHY_EDGE_ROW_163_Right_163 ();
 decap_3 PHY_EDGE_ROW_164_Right_164 ();
 decap_3 PHY_EDGE_ROW_165_Right_165 ();
 decap_3 PHY_EDGE_ROW_166_Right_166 ();
 decap_3 PHY_EDGE_ROW_167_Right_167 ();
 decap_3 PHY_EDGE_ROW_168_Right_168 ();
 decap_3 PHY_EDGE_ROW_169_Right_169 ();
 decap_3 PHY_EDGE_ROW_170_Right_170 ();
 decap_3 PHY_EDGE_ROW_171_Right_171 ();
 decap_3 PHY_EDGE_ROW_0_Left_172 ();
 decap_3 PHY_EDGE_ROW_1_Left_173 ();
 decap_3 PHY_EDGE_ROW_2_Left_174 ();
 decap_3 PHY_EDGE_ROW_3_Left_175 ();
 decap_3 PHY_EDGE_ROW_4_Left_176 ();
 decap_3 PHY_EDGE_ROW_5_Left_177 ();
 decap_3 PHY_EDGE_ROW_6_Left_178 ();
 decap_3 PHY_EDGE_ROW_7_Left_179 ();
 decap_3 PHY_EDGE_ROW_8_Left_180 ();
 decap_3 PHY_EDGE_ROW_9_Left_181 ();
 decap_3 PHY_EDGE_ROW_10_Left_182 ();
 decap_3 PHY_EDGE_ROW_11_Left_183 ();
 decap_3 PHY_EDGE_ROW_12_Left_184 ();
 decap_3 PHY_EDGE_ROW_13_Left_185 ();
 decap_3 PHY_EDGE_ROW_14_Left_186 ();
 decap_3 PHY_EDGE_ROW_15_Left_187 ();
 decap_3 PHY_EDGE_ROW_16_Left_188 ();
 decap_3 PHY_EDGE_ROW_17_Left_189 ();
 decap_3 PHY_EDGE_ROW_18_Left_190 ();
 decap_3 PHY_EDGE_ROW_19_Left_191 ();
 decap_3 PHY_EDGE_ROW_20_Left_192 ();
 decap_3 PHY_EDGE_ROW_21_Left_193 ();
 decap_3 PHY_EDGE_ROW_22_Left_194 ();
 decap_3 PHY_EDGE_ROW_23_Left_195 ();
 decap_3 PHY_EDGE_ROW_24_Left_196 ();
 decap_3 PHY_EDGE_ROW_25_Left_197 ();
 decap_3 PHY_EDGE_ROW_26_Left_198 ();
 decap_3 PHY_EDGE_ROW_27_Left_199 ();
 decap_3 PHY_EDGE_ROW_28_Left_200 ();
 decap_3 PHY_EDGE_ROW_29_Left_201 ();
 decap_3 PHY_EDGE_ROW_30_Left_202 ();
 decap_3 PHY_EDGE_ROW_31_Left_203 ();
 decap_3 PHY_EDGE_ROW_32_Left_204 ();
 decap_3 PHY_EDGE_ROW_33_Left_205 ();
 decap_3 PHY_EDGE_ROW_34_Left_206 ();
 decap_3 PHY_EDGE_ROW_35_Left_207 ();
 decap_3 PHY_EDGE_ROW_36_Left_208 ();
 decap_3 PHY_EDGE_ROW_37_Left_209 ();
 decap_3 PHY_EDGE_ROW_38_Left_210 ();
 decap_3 PHY_EDGE_ROW_39_Left_211 ();
 decap_3 PHY_EDGE_ROW_40_Left_212 ();
 decap_3 PHY_EDGE_ROW_41_Left_213 ();
 decap_3 PHY_EDGE_ROW_42_Left_214 ();
 decap_3 PHY_EDGE_ROW_43_Left_215 ();
 decap_3 PHY_EDGE_ROW_44_Left_216 ();
 decap_3 PHY_EDGE_ROW_45_Left_217 ();
 decap_3 PHY_EDGE_ROW_46_Left_218 ();
 decap_3 PHY_EDGE_ROW_47_Left_219 ();
 decap_3 PHY_EDGE_ROW_48_Left_220 ();
 decap_3 PHY_EDGE_ROW_49_Left_221 ();
 decap_3 PHY_EDGE_ROW_50_Left_222 ();
 decap_3 PHY_EDGE_ROW_51_Left_223 ();
 decap_3 PHY_EDGE_ROW_52_Left_224 ();
 decap_3 PHY_EDGE_ROW_53_Left_225 ();
 decap_3 PHY_EDGE_ROW_54_Left_226 ();
 decap_3 PHY_EDGE_ROW_55_Left_227 ();
 decap_3 PHY_EDGE_ROW_56_Left_228 ();
 decap_3 PHY_EDGE_ROW_57_Left_229 ();
 decap_3 PHY_EDGE_ROW_58_Left_230 ();
 decap_3 PHY_EDGE_ROW_59_Left_231 ();
 decap_3 PHY_EDGE_ROW_60_Left_232 ();
 decap_3 PHY_EDGE_ROW_61_Left_233 ();
 decap_3 PHY_EDGE_ROW_62_Left_234 ();
 decap_3 PHY_EDGE_ROW_63_Left_235 ();
 decap_3 PHY_EDGE_ROW_64_Left_236 ();
 decap_3 PHY_EDGE_ROW_65_Left_237 ();
 decap_3 PHY_EDGE_ROW_66_Left_238 ();
 decap_3 PHY_EDGE_ROW_67_Left_239 ();
 decap_3 PHY_EDGE_ROW_68_Left_240 ();
 decap_3 PHY_EDGE_ROW_69_Left_241 ();
 decap_3 PHY_EDGE_ROW_70_Left_242 ();
 decap_3 PHY_EDGE_ROW_71_Left_243 ();
 decap_3 PHY_EDGE_ROW_72_Left_244 ();
 decap_3 PHY_EDGE_ROW_73_Left_245 ();
 decap_3 PHY_EDGE_ROW_74_Left_246 ();
 decap_3 PHY_EDGE_ROW_75_Left_247 ();
 decap_3 PHY_EDGE_ROW_76_Left_248 ();
 decap_3 PHY_EDGE_ROW_77_Left_249 ();
 decap_3 PHY_EDGE_ROW_78_Left_250 ();
 decap_3 PHY_EDGE_ROW_79_Left_251 ();
 decap_3 PHY_EDGE_ROW_80_Left_252 ();
 decap_3 PHY_EDGE_ROW_81_Left_253 ();
 decap_3 PHY_EDGE_ROW_82_Left_254 ();
 decap_3 PHY_EDGE_ROW_83_Left_255 ();
 decap_3 PHY_EDGE_ROW_84_Left_256 ();
 decap_3 PHY_EDGE_ROW_85_Left_257 ();
 decap_3 PHY_EDGE_ROW_86_Left_258 ();
 decap_3 PHY_EDGE_ROW_87_Left_259 ();
 decap_3 PHY_EDGE_ROW_88_Left_260 ();
 decap_3 PHY_EDGE_ROW_89_Left_261 ();
 decap_3 PHY_EDGE_ROW_90_Left_262 ();
 decap_3 PHY_EDGE_ROW_91_Left_263 ();
 decap_3 PHY_EDGE_ROW_92_Left_264 ();
 decap_3 PHY_EDGE_ROW_93_Left_265 ();
 decap_3 PHY_EDGE_ROW_94_Left_266 ();
 decap_3 PHY_EDGE_ROW_95_Left_267 ();
 decap_3 PHY_EDGE_ROW_96_Left_268 ();
 decap_3 PHY_EDGE_ROW_97_Left_269 ();
 decap_3 PHY_EDGE_ROW_98_Left_270 ();
 decap_3 PHY_EDGE_ROW_99_Left_271 ();
 decap_3 PHY_EDGE_ROW_100_Left_272 ();
 decap_3 PHY_EDGE_ROW_101_Left_273 ();
 decap_3 PHY_EDGE_ROW_102_Left_274 ();
 decap_3 PHY_EDGE_ROW_103_Left_275 ();
 decap_3 PHY_EDGE_ROW_104_Left_276 ();
 decap_3 PHY_EDGE_ROW_105_Left_277 ();
 decap_3 PHY_EDGE_ROW_106_Left_278 ();
 decap_3 PHY_EDGE_ROW_107_Left_279 ();
 decap_3 PHY_EDGE_ROW_108_Left_280 ();
 decap_3 PHY_EDGE_ROW_109_Left_281 ();
 decap_3 PHY_EDGE_ROW_110_Left_282 ();
 decap_3 PHY_EDGE_ROW_111_Left_283 ();
 decap_3 PHY_EDGE_ROW_112_Left_284 ();
 decap_3 PHY_EDGE_ROW_113_Left_285 ();
 decap_3 PHY_EDGE_ROW_114_Left_286 ();
 decap_3 PHY_EDGE_ROW_115_Left_287 ();
 decap_3 PHY_EDGE_ROW_116_Left_288 ();
 decap_3 PHY_EDGE_ROW_117_Left_289 ();
 decap_3 PHY_EDGE_ROW_118_Left_290 ();
 decap_3 PHY_EDGE_ROW_119_Left_291 ();
 decap_3 PHY_EDGE_ROW_120_Left_292 ();
 decap_3 PHY_EDGE_ROW_121_Left_293 ();
 decap_3 PHY_EDGE_ROW_122_Left_294 ();
 decap_3 PHY_EDGE_ROW_123_Left_295 ();
 decap_3 PHY_EDGE_ROW_124_Left_296 ();
 decap_3 PHY_EDGE_ROW_125_Left_297 ();
 decap_3 PHY_EDGE_ROW_126_Left_298 ();
 decap_3 PHY_EDGE_ROW_127_Left_299 ();
 decap_3 PHY_EDGE_ROW_128_Left_300 ();
 decap_3 PHY_EDGE_ROW_129_Left_301 ();
 decap_3 PHY_EDGE_ROW_130_Left_302 ();
 decap_3 PHY_EDGE_ROW_131_Left_303 ();
 decap_3 PHY_EDGE_ROW_132_Left_304 ();
 decap_3 PHY_EDGE_ROW_133_Left_305 ();
 decap_3 PHY_EDGE_ROW_134_Left_306 ();
 decap_3 PHY_EDGE_ROW_135_Left_307 ();
 decap_3 PHY_EDGE_ROW_136_Left_308 ();
 decap_3 PHY_EDGE_ROW_137_Left_309 ();
 decap_3 PHY_EDGE_ROW_138_Left_310 ();
 decap_3 PHY_EDGE_ROW_139_Left_311 ();
 decap_3 PHY_EDGE_ROW_140_Left_312 ();
 decap_3 PHY_EDGE_ROW_141_Left_313 ();
 decap_3 PHY_EDGE_ROW_142_Left_314 ();
 decap_3 PHY_EDGE_ROW_143_Left_315 ();
 decap_3 PHY_EDGE_ROW_144_Left_316 ();
 decap_3 PHY_EDGE_ROW_145_Left_317 ();
 decap_3 PHY_EDGE_ROW_146_Left_318 ();
 decap_3 PHY_EDGE_ROW_147_Left_319 ();
 decap_3 PHY_EDGE_ROW_148_Left_320 ();
 decap_3 PHY_EDGE_ROW_149_Left_321 ();
 decap_3 PHY_EDGE_ROW_150_Left_322 ();
 decap_3 PHY_EDGE_ROW_151_Left_323 ();
 decap_3 PHY_EDGE_ROW_152_Left_324 ();
 decap_3 PHY_EDGE_ROW_153_Left_325 ();
 decap_3 PHY_EDGE_ROW_154_Left_326 ();
 decap_3 PHY_EDGE_ROW_155_Left_327 ();
 decap_3 PHY_EDGE_ROW_156_Left_328 ();
 decap_3 PHY_EDGE_ROW_157_Left_329 ();
 decap_3 PHY_EDGE_ROW_158_Left_330 ();
 decap_3 PHY_EDGE_ROW_159_Left_331 ();
 decap_3 PHY_EDGE_ROW_160_Left_332 ();
 decap_3 PHY_EDGE_ROW_161_Left_333 ();
 decap_3 PHY_EDGE_ROW_162_Left_334 ();
 decap_3 PHY_EDGE_ROW_163_Left_335 ();
 decap_3 PHY_EDGE_ROW_164_Left_336 ();
 decap_3 PHY_EDGE_ROW_165_Left_337 ();
 decap_3 PHY_EDGE_ROW_166_Left_338 ();
 decap_3 PHY_EDGE_ROW_167_Left_339 ();
 decap_3 PHY_EDGE_ROW_168_Left_340 ();
 decap_3 PHY_EDGE_ROW_169_Left_341 ();
 decap_3 PHY_EDGE_ROW_170_Left_342 ();
 decap_3 PHY_EDGE_ROW_171_Left_343 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_344 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_345 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_346 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_347 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_348 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_349 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_350 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_351 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_352 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_353 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_354 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_355 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_356 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_357 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_358 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_359 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_360 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_361 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_362 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_363 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_364 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_365 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_366 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_367 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_368 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_369 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_370 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_371 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_372 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_373 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_374 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_375 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_376 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_377 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_378 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_379 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_380 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_381 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_382 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_383 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_384 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_385 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_386 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_387 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_388 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_389 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_390 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_391 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_392 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_393 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_394 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_395 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_396 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_397 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_398 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_399 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_400 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_401 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_402 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_403 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_404 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_405 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_406 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_407 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_408 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_409 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_410 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_411 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_412 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_413 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_414 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_415 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_416 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_417 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_418 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_419 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_420 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_421 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_422 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_423 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_424 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_425 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_426 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_427 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_428 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_429 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_430 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_431 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_432 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_433 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_434 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_435 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_436 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_437 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_438 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_439 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_440 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_441 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_442 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_443 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_444 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_445 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_446 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_447 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_448 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_449 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_450 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_451 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_452 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_453 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_454 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_455 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_456 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_457 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_458 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_459 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_460 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_461 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_462 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_463 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_464 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_465 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_466 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_467 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_468 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_469 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_470 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_471 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_472 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_473 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_474 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_475 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_476 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_477 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_478 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_479 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_480 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_481 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_482 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_483 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_484 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_485 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_486 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_487 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_488 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_489 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_490 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_491 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_492 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_493 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_494 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_495 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_496 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_497 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_498 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_499 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_500 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_501 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_502 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_503 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_504 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_505 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_506 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_507 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_508 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_509 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_510 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_511 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_512 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_513 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_514 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_515 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_516 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_517 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_518 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_519 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_520 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_521 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_522 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_523 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_524 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_525 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_526 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_527 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_528 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_529 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_530 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_531 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_532 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_533 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_534 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_535 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_536 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_537 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_538 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_539 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_540 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_541 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_542 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_543 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_544 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_545 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_546 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_547 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_548 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_549 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_550 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_551 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_552 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_553 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_554 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_555 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_556 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_557 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_558 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_559 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_560 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_561 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_562 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_563 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_564 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_565 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_566 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_567 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_568 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_569 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_570 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_571 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_572 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_573 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_574 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_575 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_576 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_577 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_578 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_579 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_580 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_581 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_582 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_583 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_584 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_585 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_586 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_587 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_588 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_589 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_590 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_591 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_592 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_593 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_594 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_595 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_596 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_597 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_598 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_599 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_600 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_601 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_602 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_603 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_604 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_605 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_606 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_607 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_608 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_609 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_610 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_611 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_612 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_613 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_614 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_615 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_616 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_617 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_618 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_619 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_620 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_621 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_622 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_623 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_624 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_625 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_626 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_627 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_628 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_629 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_630 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_631 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_632 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_633 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_634 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_635 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_636 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_637 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_638 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_639 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_640 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_641 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_642 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_643 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_644 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_645 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_646 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_647 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_648 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_649 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_650 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_651 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_652 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_653 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_654 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_655 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_656 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_657 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_658 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_659 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_660 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_661 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_662 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_663 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_664 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_665 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_666 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_667 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_668 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_669 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_670 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_671 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_672 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_673 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_674 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_675 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_676 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_677 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_678 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_679 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_680 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_681 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_682 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_683 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_684 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_685 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_686 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_687 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_688 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_689 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_690 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_691 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_692 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_693 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_694 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_695 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_696 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_697 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_698 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_699 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_700 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_701 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_702 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_703 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_704 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_705 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_706 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_707 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_708 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_709 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_710 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_711 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_712 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_713 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_714 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_715 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_716 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_717 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_718 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_719 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_720 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_721 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_722 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_723 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_724 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_725 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_726 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_727 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_728 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_729 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_730 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_731 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_732 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_733 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_734 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_735 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_736 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_737 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_738 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_739 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_740 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_741 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_742 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_743 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_744 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_745 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_746 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_747 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_748 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_749 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_750 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_751 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_752 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_753 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_754 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_755 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_756 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_757 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_758 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_759 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_760 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_761 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_762 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_763 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_764 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_765 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_766 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_767 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_768 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_769 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_770 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_771 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_772 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_773 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_774 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_775 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_776 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_777 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_778 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_779 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_780 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_781 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_782 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_783 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_784 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_785 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_786 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_787 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_788 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_789 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_790 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_791 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_792 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_793 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_794 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_795 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_796 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_797 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_798 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_799 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_800 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_801 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_802 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_803 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_804 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_805 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_806 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_807 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_808 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_809 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_810 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_811 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_812 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_813 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_814 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_815 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_816 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_817 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_818 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_819 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_820 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_821 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_822 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_823 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_824 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_825 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_826 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_827 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_828 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_829 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_830 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_831 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_832 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_833 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_834 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_835 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_836 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_837 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_838 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_839 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_840 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_841 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_842 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_843 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_844 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_845 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_846 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_847 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_848 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_849 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_850 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_851 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_852 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_853 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_854 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_855 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_856 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_857 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_858 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_859 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_860 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_861 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_862 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_863 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_864 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_865 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_866 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_867 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_868 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_869 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_870 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_871 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_872 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_873 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_874 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_875 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_876 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_877 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_878 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_879 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_880 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_881 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_882 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_883 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_884 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_885 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_886 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_887 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_888 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_889 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_890 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_891 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_892 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_893 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_894 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_895 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_896 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_897 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_898 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_899 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_900 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_901 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_902 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_903 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_904 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_905 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_906 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_907 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_908 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_909 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_910 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_911 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_912 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_913 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_914 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_915 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_916 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_917 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_918 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_919 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_920 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_921 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_922 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_923 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_924 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_925 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_926 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_927 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_928 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_929 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_930 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_931 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_932 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_933 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_934 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_935 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_936 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_937 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_938 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_939 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_940 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_941 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_942 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_943 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_944 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_945 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_946 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_947 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_948 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_949 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_950 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_951 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_952 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_953 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_954 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_955 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_956 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_957 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_958 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_959 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_960 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_961 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_962 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_963 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_964 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_965 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_966 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_967 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_968 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_969 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_970 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_971 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_972 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_973 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_974 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_975 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_976 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_977 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_978 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_979 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_980 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_981 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_982 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_983 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_984 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_985 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_986 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_987 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_988 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_989 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_990 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_991 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_992 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_993 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_994 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_995 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_996 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_997 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_998 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_999 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1000 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1001 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1002 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1003 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1004 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1005 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1006 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1007 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1008 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1009 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1010 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1011 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1012 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1013 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1014 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1015 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1016 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1017 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1018 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1019 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1020 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1021 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1022 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1023 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1024 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1025 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1026 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1027 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1028 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1029 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1030 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1031 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1032 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1033 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1034 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1035 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1036 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1037 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1038 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1039 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1040 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1041 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1042 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1043 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1044 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1045 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1046 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1047 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1048 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1049 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1050 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1051 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1052 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1053 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1054 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1055 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1056 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1057 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1058 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1059 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1060 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1061 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1062 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1063 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1064 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1065 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1066 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1067 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1068 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1069 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1070 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1071 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1072 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1073 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1074 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1075 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1076 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1077 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1078 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1079 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1080 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1081 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1082 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1083 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1084 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1085 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1086 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1087 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1088 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1089 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1090 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1091 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1092 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1093 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1094 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1095 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1096 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1097 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1098 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1099 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1100 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1101 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1102 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1103 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1104 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1105 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1106 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1107 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1108 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1109 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1110 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1111 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1112 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1113 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1114 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1115 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1116 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1117 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1118 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1119 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1120 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1121 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1122 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1123 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1124 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1125 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1126 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1127 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1128 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1129 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1130 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1131 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1132 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1133 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1134 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1135 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1136 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1137 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1138 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1139 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1140 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1141 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1142 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1143 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1144 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1145 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1146 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1147 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1148 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1149 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1150 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1151 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1152 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1153 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1154 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1155 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1156 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1157 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1158 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1159 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1160 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1161 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1162 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1163 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1164 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1165 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1166 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1167 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1168 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1169 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1170 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1171 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1172 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1173 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1174 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1175 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1176 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1177 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1178 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1179 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1180 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1181 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1182 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1183 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1184 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1185 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1186 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1187 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1188 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1189 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1190 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1191 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1192 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1193 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1194 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1195 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1196 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1197 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1198 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1199 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1200 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1201 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1202 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1203 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1204 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1205 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1206 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1207 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1208 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1209 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1210 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1211 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1212 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1213 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1214 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1215 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1216 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1217 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1218 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1219 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1220 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1221 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1222 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1223 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1224 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1225 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1226 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1227 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1228 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1229 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1230 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1231 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1232 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1233 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1234 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1235 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1236 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1237 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1238 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1239 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1240 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1241 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1242 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1243 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1244 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1245 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1246 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1247 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1248 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1249 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1250 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1251 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1252 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1253 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1254 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1255 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1256 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1257 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1258 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1259 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1260 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1261 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1262 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1263 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1264 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1265 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1266 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1267 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1268 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1269 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1270 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1271 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1272 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1273 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1274 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1275 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1276 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1277 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1278 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1279 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1280 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1281 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1282 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1283 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1284 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1285 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1286 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1287 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1288 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1289 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1290 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1291 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1292 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1293 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1294 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1295 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1296 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1297 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1298 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1299 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1300 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1301 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1302 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1303 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1304 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1305 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1306 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1307 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1308 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1309 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1310 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1311 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1312 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1313 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1314 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1315 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1316 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1317 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1318 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1319 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1320 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1321 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1322 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1323 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1324 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1325 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1326 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1327 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1328 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1329 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1330 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1331 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1332 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1333 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1334 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1335 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1336 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1337 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1338 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1339 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1340 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1341 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1342 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1343 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1344 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1345 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1346 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1347 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1348 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1349 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1350 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1351 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1352 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1353 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1354 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1355 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1356 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1357 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1358 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1359 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1360 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1361 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1362 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1363 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1364 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1365 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1366 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1367 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1368 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1369 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1370 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1371 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1372 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1373 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1374 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1375 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1376 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1377 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1378 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1379 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1380 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1381 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1382 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1383 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1384 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1385 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1386 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1387 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1388 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1389 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1390 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1391 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1392 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1393 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1394 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1395 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1396 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1397 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1398 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1399 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1400 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1401 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1402 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1403 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1404 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1405 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1406 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1407 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1408 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1409 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1410 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1411 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1412 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1413 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1414 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1415 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1416 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1417 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1418 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1419 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1420 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1421 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1422 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1423 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1424 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1425 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1426 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1427 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1428 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1429 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1430 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1431 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1432 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1433 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1434 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1435 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1436 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1437 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1438 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1439 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1440 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1441 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1442 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1443 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1444 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1445 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1446 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1447 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1448 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1449 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1450 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1451 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1452 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1453 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1454 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1455 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1456 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1457 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1458 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1459 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1460 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1461 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1462 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1463 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1464 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1465 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1466 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1467 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1468 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1469 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1470 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1471 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1472 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1473 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1474 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1475 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1476 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1477 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1478 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1479 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1480 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1481 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1482 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1483 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1484 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1485 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1486 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1487 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1488 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1489 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1490 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1491 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1492 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1493 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1494 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1495 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1496 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1497 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1498 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1499 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1500 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1501 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1502 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1503 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1504 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1505 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1506 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1507 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1508 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1509 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1510 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1511 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1512 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1513 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1514 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1515 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1516 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1517 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1518 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1519 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1520 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1521 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1522 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1523 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1524 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1525 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1526 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1527 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1528 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1529 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1530 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1531 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1532 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1533 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1534 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1535 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1536 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1537 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1538 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1539 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1540 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1541 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1542 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1543 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1544 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1545 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1546 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1547 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1548 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1549 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1550 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1551 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1552 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1553 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1554 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1555 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1556 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1557 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1558 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1559 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1560 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1561 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1562 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1563 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1564 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1565 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1566 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1567 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1568 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1569 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1570 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1571 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1572 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1573 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1574 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1575 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1576 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1577 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1578 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1579 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1580 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1581 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1582 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1583 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1584 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1585 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1586 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1587 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1588 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1589 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1590 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1591 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1592 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1593 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1594 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1595 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1596 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1597 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1598 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1599 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1600 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1601 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1602 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1603 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1604 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1605 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1606 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1607 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1608 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1609 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1610 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1611 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1612 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1613 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1614 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1615 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1616 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1617 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1618 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1619 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1620 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1621 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1622 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1623 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1624 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1625 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1626 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1627 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1628 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1629 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1630 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1631 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1632 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1633 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1634 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1635 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1636 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1637 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1638 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1639 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1640 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1641 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1642 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1643 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1644 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1645 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1646 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1647 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1648 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1649 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1650 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1651 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1652 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1653 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1654 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1655 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1656 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1657 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1658 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1659 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1660 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1661 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1662 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1663 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1664 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1665 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1666 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1667 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1668 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1669 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1670 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1671 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1672 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1673 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1674 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1675 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1676 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1677 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1678 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1679 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1680 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1681 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1682 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1683 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1684 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1685 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1686 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1687 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1688 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1689 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1690 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1691 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1692 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1693 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1694 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1695 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1696 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1697 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1698 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1699 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1700 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1701 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1702 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1703 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1704 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1705 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1706 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1707 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1708 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1709 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1710 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1711 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1712 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1713 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1714 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1715 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1716 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1717 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1718 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1719 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1720 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1721 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1722 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1723 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1724 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1725 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1726 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1727 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1728 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1729 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1730 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1731 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1732 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1733 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1734 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1735 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1736 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1737 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1738 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1739 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1740 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1741 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1742 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1743 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1744 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1745 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1746 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1747 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1748 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1749 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1750 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1751 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1752 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1753 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1754 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1755 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1756 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1757 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1758 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1759 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1760 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1761 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1762 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1763 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1764 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1765 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1766 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1767 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1768 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1769 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1770 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1771 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1772 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1773 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1774 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1775 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1776 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1777 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1778 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1779 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1780 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1781 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1782 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1783 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1784 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1785 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1786 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1787 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1788 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1789 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1790 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1791 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1792 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1793 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1794 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1795 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1796 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1797 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1798 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1799 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1800 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1801 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1802 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1803 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1804 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1805 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1806 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1807 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1808 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1809 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1810 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1811 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1812 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1813 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1814 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1815 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1816 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1817 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1818 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1819 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1820 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1821 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1822 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1823 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1824 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1825 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1826 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1827 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1828 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1829 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1830 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1831 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1832 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1833 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1834 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1835 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1836 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1837 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1838 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1839 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1840 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1841 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1842 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1843 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1844 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1845 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1846 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1847 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1848 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1849 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1850 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1851 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1852 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1853 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1854 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1855 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1856 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1857 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1858 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1859 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1860 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1861 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1862 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1863 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1864 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1865 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1866 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1867 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1868 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1869 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1870 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1871 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1872 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1873 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1874 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1875 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1876 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1877 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1878 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1879 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1880 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1881 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1882 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1883 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1884 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1885 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1886 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1887 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1888 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1889 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1890 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1891 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1892 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1893 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1894 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1895 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1896 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1897 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1898 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1899 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1900 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1901 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1902 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1903 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1904 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1905 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1906 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1907 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1908 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1909 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1910 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1911 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1912 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1913 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1914 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1915 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1916 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1917 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1918 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1919 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1920 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1921 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1922 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1923 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1924 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1925 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1926 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1927 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1928 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1929 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1930 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1931 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1932 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1933 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1934 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1935 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1936 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1937 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1938 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1939 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1940 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1941 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1942 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1943 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1944 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1945 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1946 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1947 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1948 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1949 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1950 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1951 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1952 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1953 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1954 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1955 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1956 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1957 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1958 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1959 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1960 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1961 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1962 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1963 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1964 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1965 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1966 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1967 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1968 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1969 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1970 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1971 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1972 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1973 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1974 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1975 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1976 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1977 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1978 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1979 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1980 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1981 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1982 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1983 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1984 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1985 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1986 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1987 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1988 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1989 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1990 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1991 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1992 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1993 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1994 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1995 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1996 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1997 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1998 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1999 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2000 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2001 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2002 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2003 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2004 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2005 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2006 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2007 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2008 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2009 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2010 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2011 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2012 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2013 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2014 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2015 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2016 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2017 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2018 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2019 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2020 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2021 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2022 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2023 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2024 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2025 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2026 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2027 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2028 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2029 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2030 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2031 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2032 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2033 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2034 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2035 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2036 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2037 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2038 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2039 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2040 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2041 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2042 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2043 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2044 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2045 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2046 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2047 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2048 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2049 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2050 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2051 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2052 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2053 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2054 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2055 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2056 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2057 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2058 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2059 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2060 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2061 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2062 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2063 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2064 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2065 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2066 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2067 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2068 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2069 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2070 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2071 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2072 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2073 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2074 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2075 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2076 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2077 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2078 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2079 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2080 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2081 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2082 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2083 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2084 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2085 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2086 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2087 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2088 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2089 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2090 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2091 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2092 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2093 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2094 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2095 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2096 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2097 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2098 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2099 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2100 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2101 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2102 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2103 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2104 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2105 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2106 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2107 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2108 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2109 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2110 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2111 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2112 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2113 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2114 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2115 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2116 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2117 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2118 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2119 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2120 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2121 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2122 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2123 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2124 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2125 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2126 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2127 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2128 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2129 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2130 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2131 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2132 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2133 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2134 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2135 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2136 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2137 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2138 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2139 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2140 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2141 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2142 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2143 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2144 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2145 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2146 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2147 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2148 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2149 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2150 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2151 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2152 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2153 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2154 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2155 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2156 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2157 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2158 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2159 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2160 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2161 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2162 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2163 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2164 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2165 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2166 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2167 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2168 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2169 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2170 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2171 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2172 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2173 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2174 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2175 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2176 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2177 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2178 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2179 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2180 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2181 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2182 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2183 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2184 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2185 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2186 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2187 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2188 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2189 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2190 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2191 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2192 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2193 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2194 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2195 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2196 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2197 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2198 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2199 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2200 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2201 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2202 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2203 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2204 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2205 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2206 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2207 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2208 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2209 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2210 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2211 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2212 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2213 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2214 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2215 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2216 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2217 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2218 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2219 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2220 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2221 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2222 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2223 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2224 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2225 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2226 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2227 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2228 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2229 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2230 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2231 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2232 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2233 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2234 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2235 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2236 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2237 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2238 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2239 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2240 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2241 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2242 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2243 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2244 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2245 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2246 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2247 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2248 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2249 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2250 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2251 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2252 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2253 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2254 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2255 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2256 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2257 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2258 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2259 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2260 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2261 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2262 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2263 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2264 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2265 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2266 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2267 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2268 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2269 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2270 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2271 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2272 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2273 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2274 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2275 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2276 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2277 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2278 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2279 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2280 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2281 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2282 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2283 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2284 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2285 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2286 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2287 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2288 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2289 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2290 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2291 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2292 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2293 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2294 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2295 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2296 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2297 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2298 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2299 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2300 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2301 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2302 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2303 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2304 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2305 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2306 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2307 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2308 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2309 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2310 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2311 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2312 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2313 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2314 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2315 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2316 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2317 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2318 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2319 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2320 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2321 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2322 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2323 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2324 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2325 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2326 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2327 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2328 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2329 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2330 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2331 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2332 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2333 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2334 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2335 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2336 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2337 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2338 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2339 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2340 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2341 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2342 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2343 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2344 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2345 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2346 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2347 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2348 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2349 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2350 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2351 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2352 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2353 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2354 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2355 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2356 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2357 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2358 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2359 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2360 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2361 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2362 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2363 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2364 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2365 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2366 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2367 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2368 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2369 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2370 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2371 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2372 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2373 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2374 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2375 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2376 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2377 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2378 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2379 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2380 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2381 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2382 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2383 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2384 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2385 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2386 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2387 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2388 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2389 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2390 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2391 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2392 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2393 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2394 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2395 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2396 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2397 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2398 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2399 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2400 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2401 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2402 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2403 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2404 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2405 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2406 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2407 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2408 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2409 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2410 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2411 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2412 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2413 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2414 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2415 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2416 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2417 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2418 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2419 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2420 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2421 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2422 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2423 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2424 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2425 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2426 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2427 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2428 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2429 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2430 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2431 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2432 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2433 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2434 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2435 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2436 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2437 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2438 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2439 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2440 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2441 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2442 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2443 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2444 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2445 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2446 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2447 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2448 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2449 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2450 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2451 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2452 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2453 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2454 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2455 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2456 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2457 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2458 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2459 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2460 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2461 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2462 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2463 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2464 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2465 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2466 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2467 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2468 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2469 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2470 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2471 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2472 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2473 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2474 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2475 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2476 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2477 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2478 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2479 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2480 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2481 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2482 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2483 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2484 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2485 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2486 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2487 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2488 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2489 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2490 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2491 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2492 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2493 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2494 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2495 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2496 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2497 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2498 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2499 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2500 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2501 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2502 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2503 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2504 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2505 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2506 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2507 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2508 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2509 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2510 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2511 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2512 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2513 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2514 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2515 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2516 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2517 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2518 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2519 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2520 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2521 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2522 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2523 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2524 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2525 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2526 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2527 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2528 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2529 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2530 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2531 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2532 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2533 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2534 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2535 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2536 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2537 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2538 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2539 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2540 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2541 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2542 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2543 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2544 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2545 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2546 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2547 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2548 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2549 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2550 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2551 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2552 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2553 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2554 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2555 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2556 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2557 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2558 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2559 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2560 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2561 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2562 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2563 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2564 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2565 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2566 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2567 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2568 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2569 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2570 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2571 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2572 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2573 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2574 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2575 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2576 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2577 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2578 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2579 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2580 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2581 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2582 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2583 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2584 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2585 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2586 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2587 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2588 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2589 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2590 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2591 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2592 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2593 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2594 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2595 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2596 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2597 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2598 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2599 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2600 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2601 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2602 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2603 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2604 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2605 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2606 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2607 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2608 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2609 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2610 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2611 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2612 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2613 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2614 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2615 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2616 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2617 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2618 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2619 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2620 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2621 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2622 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2623 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2624 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2625 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2626 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2627 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2628 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2629 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2630 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2631 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2632 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2633 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2634 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2635 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2636 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2637 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2638 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2639 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2640 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2641 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2642 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2643 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2644 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2645 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2646 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2647 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2648 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2649 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2650 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2651 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2652 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2653 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2654 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2655 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2656 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2657 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2658 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2659 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2660 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2661 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2662 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2663 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2664 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2665 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2666 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2667 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2668 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2669 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2670 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2671 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2672 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2673 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2674 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2675 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2676 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2677 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2678 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2679 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2680 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2681 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2682 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2683 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2684 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2685 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2686 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2687 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2688 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2689 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2690 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2691 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2692 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2693 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2694 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2695 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2696 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2697 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2698 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2699 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2700 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2701 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2702 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2703 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2704 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2705 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2706 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2707 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2708 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2709 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2710 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2711 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2712 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2713 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2714 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2715 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2716 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2717 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2718 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2719 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2720 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2721 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2722 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2723 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2724 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2725 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2726 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2727 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2728 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2729 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2730 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2731 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2732 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2733 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2734 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2735 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2736 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2737 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2738 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2739 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2740 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2741 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2742 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2743 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2744 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2745 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2746 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2747 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2748 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2749 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2750 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2751 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2752 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2753 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2754 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2755 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2756 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2757 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2758 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2759 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2760 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2761 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2762 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2763 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2764 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2765 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2766 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2767 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2768 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2769 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2770 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2771 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2772 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2773 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2774 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2775 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2776 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2777 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2778 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2779 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2780 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2781 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2782 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2783 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2784 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2785 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2786 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2787 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2788 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2789 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2790 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2791 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2792 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2793 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2794 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2795 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2796 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2797 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2798 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2799 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2800 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2801 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2802 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2803 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2804 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2805 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2806 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2807 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2808 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2809 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2810 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2811 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2812 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2813 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2814 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2815 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2816 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2817 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2818 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2819 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2820 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2821 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2822 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2823 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2824 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2825 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2826 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2827 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2828 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2829 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2830 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2831 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2832 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2833 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2834 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2835 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2836 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2837 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2838 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2839 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2840 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2841 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2842 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2843 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2844 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2845 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2846 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2847 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2848 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2849 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2850 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2851 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2852 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2853 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2854 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2855 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2856 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2857 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2858 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2859 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2860 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2861 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2862 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2863 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2864 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2865 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2866 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2867 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2868 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2869 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2870 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2871 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2872 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2873 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2874 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2875 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2876 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2877 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2878 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2879 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2880 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2881 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2882 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2883 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2884 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2885 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2886 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2887 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2888 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2889 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2890 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2891 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2892 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2893 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2894 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2895 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2896 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2897 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2898 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2899 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2900 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2901 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2902 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2903 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2904 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2905 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2906 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2907 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2908 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2909 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2910 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2911 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2912 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2913 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2914 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2915 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2916 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2917 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2918 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2919 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2920 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2921 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2922 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2923 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2924 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2925 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2926 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2927 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2928 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2929 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2930 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2931 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2932 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2933 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2934 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2935 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2936 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2937 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2938 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2939 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2940 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2941 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2942 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2943 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2944 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2945 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2946 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2947 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2948 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2949 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2950 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2951 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2952 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2953 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2954 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2955 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2956 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2957 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2958 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2959 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2960 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2961 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2962 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2963 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2964 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2965 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2966 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2967 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2968 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2969 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2970 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2971 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2972 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2973 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2974 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2975 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2976 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2977 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2978 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2979 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2980 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2981 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2982 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2983 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2984 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2985 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2986 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2987 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2988 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2989 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2990 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2991 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2992 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2993 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2994 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2995 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2996 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2997 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2998 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2999 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3000 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3001 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3002 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3003 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3004 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3005 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3006 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3007 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3008 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3009 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3010 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3011 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3012 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3013 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3014 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3015 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3016 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3017 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3018 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3019 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3020 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3021 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3022 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3023 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3024 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3025 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3026 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3027 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3028 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3029 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3030 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3031 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3032 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3033 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3034 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3035 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3036 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3037 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3038 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3039 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3040 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3041 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3042 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3043 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3044 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3045 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3046 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3047 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3048 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3049 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3050 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3051 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3052 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3053 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3054 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3055 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3056 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3057 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3058 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3059 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3060 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3061 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3062 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3063 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3064 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3065 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3066 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3067 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3068 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3069 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3070 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3071 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3072 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3073 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3074 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3075 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3076 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3077 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3078 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3079 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3080 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3081 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3082 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3083 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3084 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3085 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3086 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3087 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3088 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3089 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3090 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3091 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3092 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3093 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3094 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3095 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3096 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3097 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3098 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3099 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3100 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3101 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3102 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3103 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3104 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3105 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3106 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3107 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3108 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3109 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3110 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3111 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3112 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3113 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3114 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3115 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3116 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3117 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3118 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3119 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3120 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3121 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3122 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3123 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3124 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3125 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3126 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3127 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3128 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3129 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3130 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3131 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3132 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3133 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3134 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3135 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3136 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3137 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3138 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3139 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3140 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3141 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3142 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3143 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3144 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3145 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3146 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3147 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3148 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3149 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3150 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3151 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3152 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3153 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3154 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3155 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3156 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3157 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3158 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3159 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3160 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3161 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3162 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3163 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3164 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3165 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3166 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3167 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3168 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3169 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3170 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3171 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3172 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3173 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3174 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3175 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3176 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3177 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3178 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3179 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3180 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3181 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3182 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3183 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3184 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3185 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3186 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3187 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3188 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3189 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3190 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3191 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3192 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3193 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3194 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3195 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3196 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3197 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3198 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3199 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3200 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3201 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3202 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3203 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3204 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3205 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3206 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3207 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3208 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3209 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3210 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3211 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3212 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3213 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3214 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3215 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3216 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3217 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3218 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3219 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3220 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3221 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3222 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3223 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3224 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3225 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3226 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3227 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3228 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3229 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3230 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3231 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3232 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3233 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3234 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3235 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3236 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3237 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3238 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3239 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3240 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3241 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3242 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3243 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3244 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3245 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3246 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3247 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3248 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3249 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3250 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3251 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3252 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3253 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3254 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3255 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3256 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3257 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3258 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3259 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3260 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3261 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3262 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3263 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3264 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3265 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3266 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3267 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3268 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3269 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3270 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3271 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3272 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3273 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3274 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3275 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3276 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3277 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3278 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3279 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3280 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3281 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3282 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3283 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3284 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3285 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3286 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3287 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3288 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3289 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3290 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3291 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3292 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3293 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3294 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3295 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3296 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3297 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3298 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3299 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3300 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3301 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3302 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3303 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3304 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3305 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3306 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3307 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3308 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3309 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3310 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3311 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3312 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3313 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3314 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3315 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3316 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3317 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3318 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3319 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3320 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3321 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3322 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3323 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3324 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3325 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3326 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3327 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3328 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3329 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3330 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3331 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3332 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3333 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3334 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3335 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3336 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3337 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3338 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3339 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3340 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3341 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3342 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3343 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3344 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3345 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3346 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3347 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3348 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3349 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3350 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3351 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3352 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3353 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3354 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3355 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3356 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3357 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3358 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3359 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3360 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3361 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3362 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3363 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3364 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3365 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3366 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3367 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3368 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3369 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3370 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3371 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3372 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3373 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3374 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3375 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3376 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3377 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3378 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3379 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3380 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3381 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3382 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3383 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3384 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3385 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3386 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3387 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3388 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3389 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3390 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3391 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3392 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3393 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3394 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3395 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3396 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3397 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3398 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3399 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3400 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3401 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3402 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3403 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3404 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3405 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3406 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3407 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3408 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3409 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3410 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3411 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3412 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3413 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3414 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3415 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3416 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3417 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3418 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3419 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3420 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3421 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3422 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3423 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3424 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3425 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3426 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3427 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3428 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3429 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3430 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3431 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3432 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3433 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3434 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3435 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3436 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3437 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3438 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3439 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3440 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3441 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3442 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3443 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3444 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3445 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3446 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3447 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3448 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3449 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3450 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3451 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3452 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3453 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3454 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3455 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3456 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3457 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3458 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3459 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3460 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3461 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3462 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3463 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3464 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3465 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3466 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3467 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3468 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3469 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3470 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3471 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3472 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3473 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3474 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3475 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3476 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3477 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3478 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3479 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3480 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3481 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3482 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3483 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3484 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3485 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3486 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3487 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3488 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3489 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3490 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3491 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3492 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3493 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3494 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3495 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3496 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3497 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3498 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3499 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3500 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3501 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3502 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3503 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3504 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3505 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3506 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3507 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3508 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3509 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3510 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3511 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3512 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3513 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3514 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3515 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3516 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3517 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3518 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3519 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3520 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3521 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3522 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3523 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3524 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3525 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3526 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3527 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3528 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3529 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3530 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3531 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3532 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3533 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3534 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3535 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3536 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3537 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3538 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3539 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3540 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3541 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3542 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3543 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3544 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3545 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3546 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3547 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3548 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3549 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3550 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3551 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3552 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3553 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3554 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3555 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3556 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3557 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3558 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3559 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3560 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3561 ();
 tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3562 ();
 clkbuf_2 input1 (.A(demod_i),
    .X(net1));
 clkbuf_1 input2 (.A(rr_data_i[0]),
    .X(net2));
 clkbuf_1 input3 (.A(rr_data_i[10]),
    .X(net3));
 clkbuf_1 input4 (.A(rr_data_i[11]),
    .X(net4));
 dlymetal6s2s_1 input5 (.A(rr_data_i[12]),
    .X(net5));
 clkbuf_1 input6 (.A(rr_data_i[13]),
    .X(net6));
 clkbuf_1 input7 (.A(rr_data_i[14]),
    .X(net7));
 clkbuf_1 input8 (.A(rr_data_i[15]),
    .X(net8));
 clkbuf_1 input9 (.A(rr_data_i[16]),
    .X(net9));
 buf_1 input10 (.A(rr_data_i[17]),
    .X(net10));
 buf_1 input11 (.A(rr_data_i[18]),
    .X(net11));
 clkbuf_1 input12 (.A(rr_data_i[19]),
    .X(net12));
 buf_1 input13 (.A(rr_data_i[1]),
    .X(net13));
 buf_1 input14 (.A(rr_data_i[20]),
    .X(net14));
 clkbuf_1 input15 (.A(rr_data_i[21]),
    .X(net15));
 buf_1 input16 (.A(rr_data_i[22]),
    .X(net16));
 clkbuf_1 input17 (.A(rr_data_i[23]),
    .X(net17));
 clkbuf_1 input18 (.A(rr_data_i[24]),
    .X(net18));
 buf_1 input19 (.A(rr_data_i[25]),
    .X(net19));
 buf_1 input20 (.A(rr_data_i[26]),
    .X(net20));
 clkbuf_1 input21 (.A(rr_data_i[27]),
    .X(net21));
 buf_1 input22 (.A(rr_data_i[28]),
    .X(net22));
 clkbuf_1 input23 (.A(rr_data_i[29]),
    .X(net23));
 buf_1 input24 (.A(rr_data_i[2]),
    .X(net24));
 clkbuf_1 input25 (.A(rr_data_i[30]),
    .X(net25));
 clkbuf_1 input26 (.A(rr_data_i[31]),
    .X(net26));
 buf_1 input27 (.A(rr_data_i[32]),
    .X(net27));
 buf_1 input28 (.A(rr_data_i[33]),
    .X(net28));
 buf_1 input29 (.A(rr_data_i[34]),
    .X(net29));
 clkbuf_1 input30 (.A(rr_data_i[35]),
    .X(net30));
 clkbuf_1 input31 (.A(rr_data_i[36]),
    .X(net31));
 clkbuf_1 input32 (.A(rr_data_i[37]),
    .X(net32));
 dlymetal6s2s_1 input33 (.A(rr_data_i[38]),
    .X(net33));
 clkbuf_1 input34 (.A(rr_data_i[39]),
    .X(net34));
 clkbuf_1 input35 (.A(rr_data_i[3]),
    .X(net35));
 clkbuf_1 input36 (.A(rr_data_i[40]),
    .X(net36));
 buf_1 input37 (.A(rr_data_i[41]),
    .X(net37));
 buf_1 input38 (.A(rr_data_i[42]),
    .X(net38));
 clkbuf_1 input39 (.A(rr_data_i[43]),
    .X(net39));
 buf_1 input40 (.A(rr_data_i[44]),
    .X(net40));
 buf_1 input41 (.A(rr_data_i[45]),
    .X(net41));
 clkbuf_1 input42 (.A(rr_data_i[46]),
    .X(net42));
 clkbuf_1 input43 (.A(rr_data_i[47]),
    .X(net43));
 buf_1 input44 (.A(rr_data_i[48]),
    .X(net44));
 clkbuf_2 input45 (.A(rr_data_i[49]),
    .X(net45));
 clkbuf_1 input46 (.A(rr_data_i[4]),
    .X(net46));
 buf_1 input47 (.A(rr_data_i[50]),
    .X(net47));
 clkbuf_1 input48 (.A(rr_data_i[51]),
    .X(net48));
 buf_1 input49 (.A(rr_data_i[52]),
    .X(net49));
 clkbuf_1 input50 (.A(rr_data_i[53]),
    .X(net50));
 buf_1 input51 (.A(rr_data_i[54]),
    .X(net51));
 clkbuf_1 input52 (.A(rr_data_i[55]),
    .X(net52));
 clkbuf_1 input53 (.A(rr_data_i[56]),
    .X(net53));
 clkbuf_2 input54 (.A(rr_data_i[57]),
    .X(net54));
 clkbuf_1 input55 (.A(rr_data_i[58]),
    .X(net55));
 clkbuf_1 input56 (.A(rr_data_i[59]),
    .X(net56));
 clkbuf_1 input57 (.A(rr_data_i[5]),
    .X(net57));
 clkbuf_2 input58 (.A(rr_data_i[60]),
    .X(net58));
 buf_1 input59 (.A(rr_data_i[61]),
    .X(net59));
 buf_1 input60 (.A(rr_data_i[62]),
    .X(net60));
 buf_1 input61 (.A(rr_data_i[63]),
    .X(net61));
 buf_1 input62 (.A(rr_data_i[6]),
    .X(net62));
 clkbuf_1 input63 (.A(rr_data_i[7]),
    .X(net63));
 clkbuf_1 input64 (.A(rr_data_i[8]),
    .X(net64));
 buf_1 input65 (.A(rr_data_i[9]),
    .X(net65));
 buf_4 input66 (.A(rst_b_i),
    .X(net66));
 clkbuf_4 input67 (.A(se_i),
    .X(net67));
 buf_4 input68 (.A(sel_nvm_i),
    .X(net68));
 clkbuf_1 input69 (.A(ti_i),
    .X(net69));
 buf_2 output70 (.A(net70),
    .X(amux_en_o));
 buf_1 output71 (.A(net71),
    .X(amux_ib_sel_o));
 buf_1 output72 (.A(net72),
    .X(amux_vcc_sel_o));
 buf_1 output73 (.A(net73),
    .X(amux_vdd_sel_o));
 buf_1 output74 (.A(net74),
    .X(amux_vref_sel_o));
 buf_2 output75 (.A(net75),
    .X(clk_trim_o[0]));
 buf_2 output76 (.A(net76),
    .X(clk_trim_o[1]));
 buf_2 output77 (.A(net77),
    .X(clk_trim_o[2]));
 buf_2 output78 (.A(net78),
    .X(demod_en_o));
 buf_1 output79 (.A(net79),
    .X(mod_o));
 buf_2 output80 (.A(net80),
    .X(rnclk_en_o));
 buf_2 output81 (.A(net81),
    .X(rnclk_trim_o[0]));
 buf_2 output82 (.A(net82),
    .X(rnclk_trim_o[1]));
 buf_2 output83 (.A(net83),
    .X(rnclk_trim_o[2]));
 buf_2 output84 (.A(net84),
    .X(rr_bank_sel_o[0]));
 buf_2 output85 (.A(net85),
    .X(rr_bank_sel_o[1]));
 buf_2 output86 (.A(net86),
    .X(rr_bank_sel_o[2]));
 buf_2 output87 (.A(net87),
    .X(rr_bank_sel_o[3]));
 buf_2 output88 (.A(net88),
    .X(rr_bl_o[0]));
 buf_2 output89 (.A(net89),
    .X(rr_bl_o[10]));
 buf_2 output90 (.A(net90),
    .X(rr_bl_o[11]));
 buf_2 output91 (.A(net91),
    .X(rr_bl_o[12]));
 buf_2 output92 (.A(net92),
    .X(rr_bl_o[13]));
 buf_2 output93 (.A(net93),
    .X(rr_bl_o[14]));
 buf_2 output94 (.A(net94),
    .X(rr_bl_o[15]));
 buf_2 output95 (.A(net95),
    .X(rr_bl_o[1]));
 buf_2 output96 (.A(net96),
    .X(rr_bl_o[2]));
 buf_2 output97 (.A(net97),
    .X(rr_bl_o[3]));
 buf_2 output98 (.A(net98),
    .X(rr_bl_o[4]));
 buf_2 output99 (.A(net99),
    .X(rr_bl_o[5]));
 buf_2 output100 (.A(net100),
    .X(rr_bl_o[6]));
 buf_2 output101 (.A(net101),
    .X(rr_bl_o[7]));
 buf_2 output102 (.A(net102),
    .X(rr_bl_o[8]));
 buf_2 output103 (.A(net103),
    .X(rr_bl_o[9]));
 buf_2 output104 (.A(net104),
    .X(rr_erase_o));
 buf_2 output105 (.A(net105),
    .X(rr_form_en_o));
 buf_2 output106 (.A(net106),
    .X(rr_prog_o));
 buf_2 output107 (.A(net107),
    .X(rr_read_o));
 buf_2 output108 (.A(net108),
    .X(rr_wl_o[0]));
 buf_2 output109 (.A(net109),
    .X(rr_wl_o[10]));
 buf_2 output110 (.A(net110),
    .X(rr_wl_o[11]));
 buf_2 output111 (.A(net111),
    .X(rr_wl_o[12]));
 buf_2 output112 (.A(net112),
    .X(rr_wl_o[13]));
 buf_2 output113 (.A(net113),
    .X(rr_wl_o[14]));
 buf_2 output114 (.A(net114),
    .X(rr_wl_o[15]));
 buf_2 output115 (.A(net115),
    .X(rr_wl_o[16]));
 buf_2 output116 (.A(net116),
    .X(rr_wl_o[17]));
 buf_2 output117 (.A(net117),
    .X(rr_wl_o[18]));
 buf_2 output118 (.A(net118),
    .X(rr_wl_o[19]));
 buf_2 output119 (.A(net119),
    .X(rr_wl_o[1]));
 buf_2 output120 (.A(net120),
    .X(rr_wl_o[20]));
 buf_2 output121 (.A(net121),
    .X(rr_wl_o[21]));
 buf_2 output122 (.A(net122),
    .X(rr_wl_o[22]));
 buf_2 output123 (.A(net123),
    .X(rr_wl_o[23]));
 buf_2 output124 (.A(net124),
    .X(rr_wl_o[24]));
 buf_2 output125 (.A(net125),
    .X(rr_wl_o[25]));
 buf_2 output126 (.A(net126),
    .X(rr_wl_o[26]));
 buf_2 output127 (.A(net127),
    .X(rr_wl_o[27]));
 buf_2 output128 (.A(net128),
    .X(rr_wl_o[28]));
 buf_2 output129 (.A(net129),
    .X(rr_wl_o[29]));
 buf_2 output130 (.A(net130),
    .X(rr_wl_o[2]));
 buf_2 output131 (.A(net131),
    .X(rr_wl_o[30]));
 buf_2 output132 (.A(net132),
    .X(rr_wl_o[31]));
 buf_2 output133 (.A(net133),
    .X(rr_wl_o[3]));
 buf_2 output134 (.A(net134),
    .X(rr_wl_o[4]));
 buf_2 output135 (.A(net135),
    .X(rr_wl_o[5]));
 buf_2 output136 (.A(net136),
    .X(rr_wl_o[6]));
 buf_2 output137 (.A(net137),
    .X(rr_wl_o[7]));
 buf_2 output138 (.A(net138),
    .X(rr_wl_o[8]));
 buf_2 output139 (.A(net139),
    .X(rr_wl_o[9]));
 buf_2 output140 (.A(net140),
    .X(to_dig_en_b_o));
 buf_1 output141 (.A(net141),
    .X(to_o));
 clkbuf_1 max_cap142 (.A(_05046_),
    .X(net142));
 clkbuf_4 fanout143 (.A(_04908_),
    .X(net143));
 clkbuf_2 fanout144 (.A(_04908_),
    .X(net144));
 buf_2 fanout145 (.A(net146),
    .X(net145));
 clkbuf_4 fanout146 (.A(_04903_),
    .X(net146));
 buf_2 fanout147 (.A(_04897_),
    .X(net147));
 clkbuf_2 fanout148 (.A(_04897_),
    .X(net148));
 buf_2 fanout149 (.A(_07955_),
    .X(net149));
 buf_2 fanout150 (.A(_07955_),
    .X(net150));
 clkbuf_4 fanout151 (.A(_07952_),
    .X(net151));
 buf_2 fanout152 (.A(_07952_),
    .X(net152));
 clkbuf_4 fanout153 (.A(_05110_),
    .X(net153));
 clkbuf_2 fanout154 (.A(_05110_),
    .X(net154));
 buf_2 fanout155 (.A(_11112_),
    .X(net155));
 buf_2 fanout156 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.fm0x_mod_en_i ),
    .X(net156));
 clkbuf_4 fanout157 (.A(_04475_),
    .X(net157));
 clkbuf_2 fanout158 (.A(_04475_),
    .X(net158));
 clkbuf_4 fanout159 (.A(_07237_),
    .X(net159));
 clkbuf_2 wire160 (.A(_02481_),
    .X(net160));
 clkbuf_4 fanout161 (.A(_11204_),
    .X(net161));
 buf_2 fanout162 (.A(net165),
    .X(net162));
 buf_2 fanout163 (.A(net165),
    .X(net163));
 clkbuf_2 fanout164 (.A(net165),
    .X(net164));
 clkbuf_2 fanout165 (.A(_11443_),
    .X(net165));
 clkbuf_4 fanout166 (.A(net169),
    .X(net166));
 buf_2 fanout167 (.A(net168),
    .X(net167));
 buf_2 fanout168 (.A(net169),
    .X(net168));
 clkbuf_2 fanout169 (.A(_11195_),
    .X(net169));
 buf_2 fanout170 (.A(net171),
    .X(net170));
 buf_2 fanout171 (.A(_06159_),
    .X(net171));
 clkbuf_4 fanout172 (.A(_11448_),
    .X(net172));
 buf_2 fanout173 (.A(_11448_),
    .X(net173));
 clkbuf_4 fanout174 (.A(net175),
    .X(net174));
 buf_4 fanout175 (.A(_11448_),
    .X(net175));
 buf_2 fanout176 (.A(net178),
    .X(net176));
 buf_2 fanout177 (.A(net178),
    .X(net177));
 clkbuf_2 fanout178 (.A(_11447_),
    .X(net178));
 clkbuf_2 fanout179 (.A(net180),
    .X(net179));
 clkbuf_4 fanout180 (.A(net181),
    .X(net180));
 clkbuf_4 fanout181 (.A(_08049_),
    .X(net181));
 clkbuf_4 fanout182 (.A(_07559_),
    .X(net182));
 clkbuf_4 fanout183 (.A(_07110_),
    .X(net183));
 buf_2 fanout184 (.A(net187),
    .X(net184));
 buf_2 fanout185 (.A(net187),
    .X(net185));
 buf_1 fanout186 (.A(net187),
    .X(net186));
 clkbuf_2 fanout187 (.A(_07109_),
    .X(net187));
 buf_2 fanout188 (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.ctr[4] ),
    .X(net188));
 clkbuf_2 fanout189 (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[2] ),
    .X(net189));
 clkbuf_2 fanout190 (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[1] ),
    .X(net190));
 clkbuf_2 fanout191 (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.state[0] ),
    .X(net191));
 buf_4 fanout192 (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.mod_en ),
    .X(net192));
 buf_2 fanout193 (.A(_08155_),
    .X(net193));
 clkbuf_4 fanout194 (.A(_02900_),
    .X(net194));
 buf_2 fanout195 (.A(_08114_),
    .X(net195));
 buf_1 fanout196 (.A(_08114_),
    .X(net196));
 buf_2 fanout197 (.A(_02949_),
    .X(net197));
 buf_2 fanout198 (.A(_02869_),
    .X(net198));
 dlymetal6s2s_1 fanout199 (.A(_02869_),
    .X(net199));
 clkbuf_4 fanout200 (.A(_11279_),
    .X(net200));
 clkbuf_4 fanout201 (.A(_07552_),
    .X(net201));
 dlymetal6s2s_1 fanout202 (.A(_07552_),
    .X(net202));
 buf_2 fanout203 (.A(net204),
    .X(net203));
 clkbuf_4 fanout204 (.A(_02922_),
    .X(net204));
 buf_4 fanout205 (.A(_02867_),
    .X(net205));
 clkbuf_2 fanout206 (.A(_02867_),
    .X(net206));
 clkbuf_8 fanout207 (.A(_02857_),
    .X(net207));
 buf_2 fanout208 (.A(_02857_),
    .X(net208));
 buf_4 fanout209 (.A(_02850_),
    .X(net209));
 buf_4 fanout210 (.A(_02849_),
    .X(net210));
 buf_2 fanout211 (.A(net212),
    .X(net211));
 buf_2 fanout212 (.A(net216),
    .X(net212));
 buf_2 fanout213 (.A(net215),
    .X(net213));
 clkbuf_4 fanout214 (.A(net215),
    .X(net214));
 clkbuf_2 fanout215 (.A(net216),
    .X(net215));
 dlymetal6s2s_1 fanout216 (.A(_02842_),
    .X(net216));
 buf_2 fanout217 (.A(_02841_),
    .X(net217));
 clkbuf_4 fanout218 (.A(_02841_),
    .X(net218));
 buf_2 fanout219 (.A(net221),
    .X(net219));
 clkbuf_2 fanout220 (.A(net221),
    .X(net220));
 clkbuf_4 fanout221 (.A(_02841_),
    .X(net221));
 buf_2 fanout222 (.A(net224),
    .X(net222));
 clkbuf_2 fanout223 (.A(net224),
    .X(net223));
 buf_2 fanout224 (.A(_11274_),
    .X(net224));
 buf_2 fanout225 (.A(_11274_),
    .X(net225));
 clkbuf_2 fanout226 (.A(_11274_),
    .X(net226));
 buf_2 fanout227 (.A(net234),
    .X(net227));
 clkbuf_2 fanout228 (.A(net234),
    .X(net228));
 buf_2 fanout229 (.A(net234),
    .X(net229));
 dlymetal6s2s_1 fanout230 (.A(net234),
    .X(net230));
 buf_2 fanout231 (.A(net234),
    .X(net231));
 clkbuf_2 fanout232 (.A(net234),
    .X(net232));
 buf_2 fanout233 (.A(net234),
    .X(net233));
 clkbuf_2 fanout234 (.A(_11273_),
    .X(net234));
 buf_4 fanout235 (.A(net236),
    .X(net235));
 clkbuf_4 fanout236 (.A(_11250_),
    .X(net236));
 buf_2 fanout237 (.A(net239),
    .X(net237));
 clkbuf_4 fanout238 (.A(net239),
    .X(net238));
 buf_2 fanout239 (.A(_11235_),
    .X(net239));
 buf_2 fanout240 (.A(net241),
    .X(net240));
 buf_2 fanout241 (.A(_11235_),
    .X(net241));
 buf_2 fanout242 (.A(net244),
    .X(net242));
 dlymetal6s2s_1 fanout243 (.A(net244),
    .X(net243));
 buf_2 fanout244 (.A(net247),
    .X(net244));
 clkbuf_4 fanout245 (.A(net247),
    .X(net245));
 clkbuf_4 fanout246 (.A(net247),
    .X(net246));
 buf_2 fanout247 (.A(_11234_),
    .X(net247));
 clkbuf_4 fanout248 (.A(net250),
    .X(net248));
 buf_2 fanout249 (.A(net250),
    .X(net249));
 dlymetal6s2s_1 fanout250 (.A(_11227_),
    .X(net250));
 buf_2 fanout251 (.A(net253),
    .X(net251));
 buf_2 fanout252 (.A(net253),
    .X(net252));
 clkbuf_2 fanout253 (.A(_11226_),
    .X(net253));
 buf_2 fanout254 (.A(net255),
    .X(net254));
 clkbuf_2 fanout255 (.A(_06306_),
    .X(net255));
 clkbuf_4 fanout256 (.A(_02947_),
    .X(net256));
 clkbuf_2 fanout257 (.A(_02947_),
    .X(net257));
 buf_2 fanout258 (.A(_02946_),
    .X(net258));
 buf_2 fanout259 (.A(net261),
    .X(net259));
 clkbuf_2 fanout260 (.A(net261),
    .X(net260));
 buf_2 fanout261 (.A(net264),
    .X(net261));
 buf_2 fanout262 (.A(net263),
    .X(net262));
 buf_2 fanout263 (.A(net264),
    .X(net263));
 dlymetal6s2s_1 fanout264 (.A(_02892_),
    .X(net264));
 buf_2 fanout265 (.A(net268),
    .X(net265));
 clkbuf_2 fanout266 (.A(net268),
    .X(net266));
 buf_2 fanout267 (.A(net268),
    .X(net267));
 dlymetal6s2s_1 fanout268 (.A(_02891_),
    .X(net268));
 buf_2 fanout269 (.A(net270),
    .X(net269));
 clkbuf_2 fanout270 (.A(_02891_),
    .X(net270));
 buf_2 fanout271 (.A(_02891_),
    .X(net271));
 clkbuf_2 fanout272 (.A(_02891_),
    .X(net272));
 buf_2 fanout273 (.A(net276),
    .X(net273));
 dlymetal6s2s_1 fanout274 (.A(net276),
    .X(net274));
 buf_2 fanout275 (.A(net276),
    .X(net275));
 clkbuf_2 fanout276 (.A(_02834_),
    .X(net276));
 clkbuf_4 fanout277 (.A(_02833_),
    .X(net277));
 buf_2 fanout278 (.A(net279),
    .X(net278));
 buf_2 fanout279 (.A(_02833_),
    .X(net279));
 buf_2 fanout280 (.A(_11358_),
    .X(net280));
 clkbuf_2 fanout281 (.A(_11358_),
    .X(net281));
 buf_2 fanout282 (.A(_11306_),
    .X(net282));
 buf_2 fanout283 (.A(_11306_),
    .X(net283));
 buf_2 fanout284 (.A(net286),
    .X(net284));
 buf_2 fanout285 (.A(net286),
    .X(net285));
 clkbuf_2 fanout286 (.A(_11305_),
    .X(net286));
 buf_4 fanout287 (.A(_11259_),
    .X(net287));
 buf_4 fanout288 (.A(_11243_),
    .X(net288));
 buf_4 fanout289 (.A(_11242_),
    .X(net289));
 clkbuf_2 fanout290 (.A(_06305_),
    .X(net290));
 buf_1 fanout291 (.A(_06305_),
    .X(net291));
 buf_2 fanout292 (.A(net293),
    .X(net292));
 clkbuf_2 fanout293 (.A(net294),
    .X(net293));
 clkbuf_2 fanout294 (.A(net296),
    .X(net294));
 buf_2 fanout295 (.A(net296),
    .X(net295));
 buf_2 fanout296 (.A(_05704_),
    .X(net296));
 buf_2 fanout297 (.A(net300),
    .X(net297));
 clkbuf_2 fanout298 (.A(net300),
    .X(net298));
 clkbuf_4 fanout299 (.A(net300),
    .X(net299));
 buf_2 fanout300 (.A(_05671_),
    .X(net300));
 buf_4 fanout301 (.A(_05437_),
    .X(net301));
 buf_2 fanout302 (.A(_05437_),
    .X(net302));
 buf_4 fanout303 (.A(_05436_),
    .X(net303));
 buf_2 fanout304 (.A(_05436_),
    .X(net304));
 clkbuf_4 fanout305 (.A(net307),
    .X(net305));
 buf_2 fanout306 (.A(net308),
    .X(net306));
 dlymetal6s2s_1 fanout307 (.A(net308),
    .X(net307));
 buf_4 fanout308 (.A(_05835_),
    .X(net308));
 buf_4 fanout309 (.A(_05788_),
    .X(net309));
 buf_2 fanout310 (.A(_05788_),
    .X(net310));
 clkbuf_4 fanout311 (.A(net313),
    .X(net311));
 clkbuf_4 fanout312 (.A(net313),
    .X(net312));
 buf_4 fanout313 (.A(_05737_),
    .X(net313));
 clkbuf_8 fanout314 (.A(_05622_),
    .X(net314));
 buf_2 fanout315 (.A(_05622_),
    .X(net315));
 clkbuf_8 fanout316 (.A(_05621_),
    .X(net316));
 buf_2 fanout317 (.A(_05621_),
    .X(net317));
 buf_4 fanout318 (.A(_05572_),
    .X(net318));
 buf_2 fanout319 (.A(_05572_),
    .X(net319));
 buf_4 fanout320 (.A(_05571_),
    .X(net320));
 buf_2 fanout321 (.A(_05571_),
    .X(net321));
 buf_2 fanout322 (.A(net325),
    .X(net322));
 buf_2 fanout323 (.A(net324),
    .X(net323));
 buf_2 fanout324 (.A(net325),
    .X(net324));
 clkbuf_2 fanout325 (.A(net328),
    .X(net325));
 buf_2 fanout326 (.A(net327),
    .X(net326));
 buf_2 fanout327 (.A(net328),
    .X(net327));
 dlymetal6s2s_1 fanout328 (.A(_04446_),
    .X(net328));
 buf_2 fanout329 (.A(_04446_),
    .X(net329));
 buf_2 fanout330 (.A(_04446_),
    .X(net330));
 buf_2 fanout331 (.A(net333),
    .X(net331));
 clkbuf_2 fanout332 (.A(net333),
    .X(net332));
 buf_2 fanout333 (.A(_04446_),
    .X(net333));
 clkbuf_2 wire334 (.A(_02734_),
    .X(net334));
 buf_1 max_cap335 (.A(_10789_),
    .X(net335));
 buf_2 fanout336 (.A(_08549_),
    .X(net336));
 clkbuf_2 fanout337 (.A(_08549_),
    .X(net337));
 clkbuf_4 fanout338 (.A(_08136_),
    .X(net338));
 buf_2 fanout339 (.A(_08134_),
    .X(net339));
 clkbuf_2 fanout340 (.A(_08134_),
    .X(net340));
 buf_2 fanout341 (.A(_08125_),
    .X(net341));
 buf_2 fanout342 (.A(_08122_),
    .X(net342));
 clkbuf_4 fanout343 (.A(net346),
    .X(net343));
 clkbuf_2 fanout344 (.A(net346),
    .X(net344));
 clkbuf_4 fanout345 (.A(net346),
    .X(net345));
 buf_2 fanout346 (.A(_05434_),
    .X(net346));
 buf_2 fanout347 (.A(net348),
    .X(net347));
 buf_2 fanout348 (.A(net349),
    .X(net348));
 clkbuf_2 fanout349 (.A(_11442_),
    .X(net349));
 clkbuf_4 fanout350 (.A(net351),
    .X(net350));
 buf_1 fanout351 (.A(net352),
    .X(net351));
 buf_2 fanout352 (.A(net353),
    .X(net352));
 clkbuf_4 fanout353 (.A(_11224_),
    .X(net353));
 buf_2 fanout354 (.A(net355),
    .X(net354));
 buf_2 fanout355 (.A(_11217_),
    .X(net355));
 buf_2 fanout356 (.A(_11213_),
    .X(net356));
 clkbuf_2 fanout357 (.A(_11213_),
    .X(net357));
 buf_4 fanout358 (.A(net359),
    .X(net358));
 clkbuf_4 fanout359 (.A(_11206_),
    .X(net359));
 clkbuf_4 fanout360 (.A(net362),
    .X(net360));
 buf_2 fanout361 (.A(net362),
    .X(net361));
 buf_2 fanout362 (.A(net363),
    .X(net362));
 buf_4 fanout363 (.A(_11205_),
    .X(net363));
 buf_2 fanout364 (.A(_11200_),
    .X(net364));
 buf_2 fanout365 (.A(_11200_),
    .X(net365));
 buf_4 fanout366 (.A(_07523_),
    .X(net366));
 clkbuf_2 fanout367 (.A(net368),
    .X(net367));
 dlymetal6s2s_1 fanout368 (.A(net371),
    .X(net368));
 buf_2 fanout369 (.A(net370),
    .X(net369));
 buf_2 fanout370 (.A(net371),
    .X(net370));
 buf_1 fanout371 (.A(net374),
    .X(net371));
 buf_2 fanout372 (.A(net373),
    .X(net372));
 clkbuf_4 fanout373 (.A(net374),
    .X(net373));
 clkbuf_2 fanout374 (.A(_07522_),
    .X(net374));
 clkbuf_2 fanout375 (.A(net376),
    .X(net375));
 clkbuf_2 fanout376 (.A(net381),
    .X(net376));
 buf_2 fanout377 (.A(net378),
    .X(net377));
 buf_2 fanout378 (.A(net381),
    .X(net378));
 buf_2 fanout379 (.A(net381),
    .X(net379));
 clkbuf_2 fanout380 (.A(net381),
    .X(net380));
 clkbuf_2 fanout381 (.A(net387),
    .X(net381));
 clkbuf_2 fanout382 (.A(net383),
    .X(net382));
 clkbuf_2 fanout383 (.A(net384),
    .X(net383));
 clkbuf_2 fanout384 (.A(net387),
    .X(net384));
 buf_2 fanout385 (.A(net386),
    .X(net385));
 dlymetal6s2s_1 fanout386 (.A(net387),
    .X(net386));
 clkbuf_2 fanout387 (.A(_07522_),
    .X(net387));
 buf_2 fanout388 (.A(_11215_),
    .X(net388));
 buf_2 fanout389 (.A(_11215_),
    .X(net389));
 buf_2 fanout390 (.A(net391),
    .X(net390));
 buf_2 fanout391 (.A(_11211_),
    .X(net391));
 buf_2 fanout392 (.A(net393),
    .X(net392));
 clkbuf_4 fanout393 (.A(net394),
    .X(net393));
 buf_2 fanout394 (.A(_11208_),
    .X(net394));
 clkbuf_4 fanout395 (.A(_11207_),
    .X(net395));
 clkbuf_4 fanout396 (.A(_11207_),
    .X(net396));
 buf_4 fanout397 (.A(_11207_),
    .X(net397));
 buf_2 fanout398 (.A(_07519_),
    .X(net398));
 buf_2 fanout399 (.A(net400),
    .X(net399));
 buf_1 fanout400 (.A(net401),
    .X(net400));
 clkbuf_4 fanout401 (.A(net402),
    .X(net401));
 clkbuf_4 fanout402 (.A(_11222_),
    .X(net402));
 buf_2 fanout403 (.A(_11201_),
    .X(net403));
 clkbuf_2 fanout404 (.A(_11201_),
    .X(net404));
 clkbuf_4 fanout405 (.A(_07094_),
    .X(net405));
 buf_2 fanout406 (.A(_07094_),
    .X(net406));
 buf_2 fanout407 (.A(net409),
    .X(net407));
 buf_2 fanout408 (.A(net409),
    .X(net408));
 clkbuf_4 fanout409 (.A(_07094_),
    .X(net409));
 clkbuf_4 fanout410 (.A(net412),
    .X(net410));
 clkbuf_2 fanout411 (.A(net412),
    .X(net411));
 clkbuf_4 fanout412 (.A(_07094_),
    .X(net412));
 buf_2 fanout413 (.A(\digitop_pav2.aes128_inst.aes128_counter.cnt_fin_3b_o ),
    .X(net413));
 buf_2 fanout414 (.A(net415),
    .X(net414));
 buf_2 fanout415 (.A(net417),
    .X(net415));
 clkbuf_4 fanout416 (.A(net417),
    .X(net416));
 buf_2 fanout417 (.A(net428),
    .X(net417));
 buf_2 fanout418 (.A(net420),
    .X(net418));
 buf_2 fanout419 (.A(net420),
    .X(net419));
 buf_2 fanout420 (.A(net424),
    .X(net420));
 buf_2 fanout421 (.A(net424),
    .X(net421));
 buf_2 fanout422 (.A(net424),
    .X(net422));
 buf_2 fanout423 (.A(net424),
    .X(net423));
 clkbuf_2 fanout424 (.A(net428),
    .X(net424));
 buf_2 fanout425 (.A(net427),
    .X(net425));
 buf_2 fanout426 (.A(net427),
    .X(net426));
 clkbuf_2 fanout427 (.A(net428),
    .X(net427));
 buf_2 fanout428 (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[7] ),
    .X(net428));
 buf_2 fanout429 (.A(net430),
    .X(net429));
 buf_2 fanout430 (.A(net431),
    .X(net430));
 buf_2 fanout431 (.A(net441),
    .X(net431));
 buf_2 fanout432 (.A(net434),
    .X(net432));
 buf_2 fanout433 (.A(net434),
    .X(net433));
 clkbuf_2 fanout434 (.A(net435),
    .X(net434));
 buf_2 fanout435 (.A(net441),
    .X(net435));
 buf_2 fanout436 (.A(net441),
    .X(net436));
 buf_2 fanout437 (.A(net441),
    .X(net437));
 buf_2 fanout438 (.A(net439),
    .X(net438));
 clkbuf_4 fanout439 (.A(net440),
    .X(net439));
 buf_2 fanout440 (.A(net441),
    .X(net440));
 buf_2 fanout441 (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[6] ),
    .X(net441));
 buf_2 fanout442 (.A(net443),
    .X(net442));
 buf_2 fanout443 (.A(net459),
    .X(net443));
 clkbuf_4 fanout444 (.A(net445),
    .X(net444));
 clkbuf_2 fanout445 (.A(net446),
    .X(net445));
 clkbuf_2 fanout446 (.A(net459),
    .X(net446));
 buf_2 fanout447 (.A(net448),
    .X(net447));
 buf_2 fanout448 (.A(net449),
    .X(net448));
 clkbuf_2 fanout449 (.A(net459),
    .X(net449));
 clkbuf_4 fanout450 (.A(net451),
    .X(net450));
 buf_2 fanout451 (.A(net459),
    .X(net451));
 clkbuf_4 fanout452 (.A(net454),
    .X(net452));
 dlymetal6s2s_1 fanout453 (.A(net454),
    .X(net453));
 buf_2 fanout454 (.A(net459),
    .X(net454));
 buf_2 fanout455 (.A(net456),
    .X(net455));
 dlymetal6s2s_1 fanout456 (.A(net458),
    .X(net456));
 clkbuf_4 fanout457 (.A(net458),
    .X(net457));
 buf_2 fanout458 (.A(net459),
    .X(net458));
 clkbuf_4 fanout459 (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[5] ),
    .X(net459));
 buf_2 fanout460 (.A(net462),
    .X(net460));
 clkbuf_4 fanout461 (.A(net462),
    .X(net461));
 clkbuf_4 fanout462 (.A(net464),
    .X(net462));
 clkbuf_4 fanout463 (.A(net464),
    .X(net463));
 clkbuf_2 fanout464 (.A(net465),
    .X(net464));
 buf_4 fanout465 (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[5] ),
    .X(net465));
 buf_2 fanout466 (.A(net470),
    .X(net466));
 buf_2 fanout467 (.A(net470),
    .X(net467));
 buf_4 fanout468 (.A(net470),
    .X(net468));
 clkbuf_2 fanout469 (.A(net470),
    .X(net469));
 clkbuf_4 fanout470 (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[3] ),
    .X(net470));
 buf_4 fanout471 (.A(net473),
    .X(net471));
 clkbuf_2 fanout472 (.A(net473),
    .X(net472));
 clkbuf_4 fanout473 (.A(\digitop_pav2.aes128_inst.aes128_regs.state_areg_r[1] ),
    .X(net473));
 clkbuf_1 max_cap474 (.A(_10176_),
    .X(net474));
 clkbuf_4 fanout475 (.A(_00991_),
    .X(net475));
 buf_2 fanout476 (.A(_09756_),
    .X(net476));
 clkbuf_2 fanout477 (.A(_09756_),
    .X(net477));
 clkbuf_4 fanout478 (.A(_09726_),
    .X(net478));
 buf_2 fanout479 (.A(_09792_),
    .X(net479));
 dlymetal6s2s_1 fanout480 (.A(_09792_),
    .X(net480));
 buf_2 fanout481 (.A(_09786_),
    .X(net481));
 buf_2 fanout482 (.A(_09777_),
    .X(net482));
 buf_2 fanout483 (.A(_09777_),
    .X(net483));
 buf_2 fanout484 (.A(_09769_),
    .X(net484));
 buf_2 fanout485 (.A(_09762_),
    .X(net485));
 dlymetal6s2s_1 fanout486 (.A(_09762_),
    .X(net486));
 clkbuf_2 fanout487 (.A(net488),
    .X(net487));
 buf_2 fanout488 (.A(net489),
    .X(net488));
 buf_2 fanout489 (.A(net490),
    .X(net489));
 clkbuf_4 fanout490 (.A(_09752_),
    .X(net490));
 buf_2 fanout491 (.A(_09649_),
    .X(net491));
 clkbuf_2 fanout492 (.A(_09798_),
    .X(net492));
 buf_2 fanout493 (.A(_09587_),
    .X(net493));
 buf_2 fanout494 (.A(_09581_),
    .X(net494));
 buf_2 fanout495 (.A(_09589_),
    .X(net495));
 buf_2 fanout496 (.A(net498),
    .X(net496));
 buf_2 fanout497 (.A(net498),
    .X(net497));
 buf_2 fanout498 (.A(_09270_),
    .X(net498));
 clkbuf_4 fanout499 (.A(_09269_),
    .X(net499));
 buf_2 fanout500 (.A(_09269_),
    .X(net500));
 clkbuf_4 fanout501 (.A(net502),
    .X(net501));
 clkbuf_2 fanout502 (.A(_09259_),
    .X(net502));
 clkbuf_2 max_cap503 (.A(_09250_),
    .X(net503));
 buf_2 fanout504 (.A(net505),
    .X(net504));
 buf_2 fanout505 (.A(_09249_),
    .X(net505));
 buf_2 fanout506 (.A(_09249_),
    .X(net506));
 dlymetal6s2s_1 fanout507 (.A(_09249_),
    .X(net507));
 clkbuf_4 fanout508 (.A(net509),
    .X(net508));
 clkbuf_4 fanout509 (.A(_09263_),
    .X(net509));
 clkbuf_4 fanout510 (.A(net511),
    .X(net510));
 clkbuf_4 fanout511 (.A(_09258_),
    .X(net511));
 clkbuf_4 fanout512 (.A(net513),
    .X(net512));
 clkbuf_4 fanout513 (.A(_09673_),
    .X(net513));
 clkbuf_2 max_cap514 (.A(_09672_),
    .X(net514));
 buf_2 fanout515 (.A(_09280_),
    .X(net515));
 clkbuf_2 fanout516 (.A(_09280_),
    .X(net516));
 buf_2 fanout517 (.A(net518),
    .X(net517));
 clkbuf_4 fanout518 (.A(net519),
    .X(net518));
 buf_2 fanout519 (.A(_09279_),
    .X(net519));
 clkbuf_4 fanout520 (.A(_09277_),
    .X(net520));
 dlymetal6s2s_1 fanout521 (.A(_09277_),
    .X(net521));
 clkbuf_4 fanout522 (.A(_09228_),
    .X(net522));
 buf_2 fanout523 (.A(_09228_),
    .X(net523));
 clkbuf_4 fanout524 (.A(net525),
    .X(net524));
 buf_2 fanout525 (.A(_08521_),
    .X(net525));
 clkbuf_4 fanout526 (.A(_05085_),
    .X(net526));
 buf_2 fanout527 (.A(_04655_),
    .X(net527));
 clkbuf_2 fanout528 (.A(_04655_),
    .X(net528));
 buf_2 fanout529 (.A(net530),
    .X(net529));
 buf_2 fanout530 (.A(_09541_),
    .X(net530));
 buf_2 fanout531 (.A(_09540_),
    .X(net531));
 buf_2 fanout532 (.A(_09540_),
    .X(net532));
 clkbuf_4 fanout533 (.A(_09187_),
    .X(net533));
 buf_2 fanout534 (.A(_11395_),
    .X(net534));
 clkbuf_2 fanout535 (.A(_11395_),
    .X(net535));
 clkbuf_8 fanout536 (.A(_09179_),
    .X(net536));
 buf_2 fanout537 (.A(_08566_),
    .X(net537));
 buf_2 fanout538 (.A(_08566_),
    .X(net538));
 buf_2 fanout539 (.A(_08562_),
    .X(net539));
 clkbuf_2 fanout540 (.A(_08562_),
    .X(net540));
 buf_2 fanout541 (.A(_08556_),
    .X(net541));
 clkbuf_2 fanout542 (.A(_08556_),
    .X(net542));
 buf_2 fanout543 (.A(_08555_),
    .X(net543));
 buf_2 fanout544 (.A(_08553_),
    .X(net544));
 clkbuf_2 fanout545 (.A(_08553_),
    .X(net545));
 buf_2 fanout546 (.A(_08552_),
    .X(net546));
 buf_2 fanout547 (.A(_08551_),
    .X(net547));
 dlymetal6s2s_1 fanout548 (.A(_08551_),
    .X(net548));
 buf_2 fanout549 (.A(_08550_),
    .X(net549));
 dlymetal6s2s_1 fanout550 (.A(_08550_),
    .X(net550));
 buf_2 fanout551 (.A(_08548_),
    .X(net551));
 clkbuf_2 fanout552 (.A(_08548_),
    .X(net552));
 buf_2 fanout553 (.A(_08547_),
    .X(net553));
 dlymetal6s2s_1 fanout554 (.A(_08547_),
    .X(net554));
 buf_2 fanout555 (.A(_08546_),
    .X(net555));
 clkbuf_4 fanout556 (.A(_08542_),
    .X(net556));
 clkbuf_2 fanout557 (.A(_08542_),
    .X(net557));
 clkbuf_4 fanout558 (.A(_08538_),
    .X(net558));
 clkbuf_2 fanout559 (.A(_08538_),
    .X(net559));
 buf_4 fanout560 (.A(_08533_),
    .X(net560));
 clkbuf_2 fanout561 (.A(_08533_),
    .X(net561));
 buf_4 fanout562 (.A(_08531_),
    .X(net562));
 clkbuf_2 fanout563 (.A(_08531_),
    .X(net563));
 buf_4 fanout564 (.A(_08530_),
    .X(net564));
 clkbuf_2 fanout565 (.A(_08530_),
    .X(net565));
 clkbuf_4 fanout566 (.A(_08529_),
    .X(net566));
 clkbuf_2 fanout567 (.A(_08529_),
    .X(net567));
 clkbuf_4 fanout568 (.A(_08527_),
    .X(net568));
 clkbuf_2 fanout569 (.A(_08527_),
    .X(net569));
 buf_2 fanout570 (.A(_06326_),
    .X(net570));
 buf_2 fanout571 (.A(_06304_),
    .X(net571));
 clkbuf_4 fanout572 (.A(net573),
    .X(net572));
 buf_2 fanout573 (.A(_04427_),
    .X(net573));
 clkbuf_4 fanout574 (.A(_11434_),
    .X(net574));
 clkbuf_4 fanout575 (.A(_11430_),
    .X(net575));
 clkbuf_2 fanout576 (.A(_11430_),
    .X(net576));
 clkbuf_4 fanout577 (.A(_11401_),
    .X(net577));
 buf_4 fanout578 (.A(_09172_),
    .X(net578));
 clkbuf_4 fanout579 (.A(_09172_),
    .X(net579));
 clkbuf_2 fanout580 (.A(net581),
    .X(net580));
 clkbuf_2 fanout581 (.A(_08545_),
    .X(net581));
 clkbuf_2 fanout582 (.A(net583),
    .X(net582));
 buf_1 max_cap583 (.A(_08525_),
    .X(net583));
 clkbuf_4 fanout584 (.A(net585),
    .X(net584));
 buf_2 fanout585 (.A(_04426_),
    .X(net585));
 clkbuf_4 fanout586 (.A(net587),
    .X(net586));
 buf_2 fanout587 (.A(_04425_),
    .X(net587));
 clkbuf_4 fanout588 (.A(_04424_),
    .X(net588));
 buf_2 fanout589 (.A(_04424_),
    .X(net589));
 clkbuf_4 fanout590 (.A(_03018_),
    .X(net590));
 buf_2 fanout591 (.A(_03013_),
    .X(net591));
 buf_2 fanout592 (.A(_03010_),
    .X(net592));
 clkbuf_4 fanout593 (.A(_03006_),
    .X(net593));
 buf_2 fanout594 (.A(_11420_),
    .X(net594));
 clkbuf_4 fanout595 (.A(_11415_),
    .X(net595));
 clkbuf_2 fanout596 (.A(_11415_),
    .X(net596));
 buf_2 fanout597 (.A(_11414_),
    .X(net597));
 clkbuf_4 fanout598 (.A(_11414_),
    .X(net598));
 buf_2 fanout599 (.A(_11411_),
    .X(net599));
 buf_2 fanout600 (.A(net601),
    .X(net600));
 clkbuf_2 fanout601 (.A(_10418_),
    .X(net601));
 buf_2 fanout602 (.A(_10417_),
    .X(net602));
 buf_1 fanout603 (.A(_10417_),
    .X(net603));
 clkbuf_2 fanout604 (.A(net608),
    .X(net604));
 clkbuf_2 fanout605 (.A(net608),
    .X(net605));
 clkbuf_2 fanout606 (.A(net607),
    .X(net606));
 dlymetal6s2s_1 fanout607 (.A(net608),
    .X(net607));
 clkbuf_2 fanout608 (.A(_06408_),
    .X(net608));
 clkbuf_2 fanout609 (.A(net610),
    .X(net609));
 clkbuf_2 fanout610 (.A(net611),
    .X(net610));
 clkbuf_2 fanout611 (.A(net613),
    .X(net611));
 buf_2 fanout612 (.A(net613),
    .X(net612));
 clkbuf_2 fanout613 (.A(_06408_),
    .X(net613));
 clkbuf_2 fanout614 (.A(net639),
    .X(net614));
 clkbuf_2 fanout615 (.A(net639),
    .X(net615));
 clkbuf_2 fanout616 (.A(net617),
    .X(net616));
 clkbuf_2 fanout617 (.A(net639),
    .X(net617));
 clkbuf_2 fanout618 (.A(net619),
    .X(net618));
 buf_1 fanout619 (.A(net624),
    .X(net619));
 clkbuf_2 fanout620 (.A(net624),
    .X(net620));
 clkbuf_2 fanout621 (.A(net623),
    .X(net621));
 clkbuf_2 fanout622 (.A(net623),
    .X(net622));
 clkbuf_2 fanout623 (.A(net624),
    .X(net623));
 clkbuf_2 fanout624 (.A(net639),
    .X(net624));
 clkbuf_2 fanout625 (.A(net638),
    .X(net625));
 buf_2 fanout626 (.A(net638),
    .X(net626));
 clkbuf_2 fanout627 (.A(net629),
    .X(net627));
 buf_1 fanout628 (.A(net629),
    .X(net628));
 clkbuf_2 fanout629 (.A(net638),
    .X(net629));
 clkbuf_2 fanout630 (.A(net633),
    .X(net630));
 clkbuf_2 fanout631 (.A(net632),
    .X(net631));
 buf_1 fanout632 (.A(net633),
    .X(net632));
 dlymetal6s2s_1 fanout633 (.A(net638),
    .X(net633));
 clkbuf_2 fanout634 (.A(net635),
    .X(net634));
 dlymetal6s2s_1 fanout635 (.A(net637),
    .X(net635));
 clkbuf_2 fanout636 (.A(net637),
    .X(net636));
 clkbuf_2 fanout637 (.A(net638),
    .X(net637));
 buf_2 fanout638 (.A(net639),
    .X(net638));
 buf_2 fanout639 (.A(_06408_),
    .X(net639));
 clkbuf_2 fanout640 (.A(net642),
    .X(net640));
 clkbuf_2 fanout641 (.A(net642),
    .X(net641));
 buf_2 fanout642 (.A(net647),
    .X(net642));
 clkbuf_2 fanout643 (.A(net644),
    .X(net643));
 buf_2 fanout644 (.A(net647),
    .X(net644));
 clkbuf_2 fanout645 (.A(net646),
    .X(net645));
 clkbuf_2 fanout646 (.A(net647),
    .X(net646));
 buf_2 fanout647 (.A(net648),
    .X(net647));
 buf_2 fanout648 (.A(_06407_),
    .X(net648));
 clkbuf_2 fanout649 (.A(net654),
    .X(net649));
 clkbuf_2 fanout650 (.A(net651),
    .X(net650));
 dlymetal6s2s_1 fanout651 (.A(net654),
    .X(net651));
 clkbuf_2 fanout652 (.A(net654),
    .X(net652));
 buf_1 fanout653 (.A(net654),
    .X(net653));
 clkbuf_2 fanout654 (.A(net662),
    .X(net654));
 clkbuf_2 fanout655 (.A(net656),
    .X(net655));
 clkbuf_2 fanout656 (.A(net662),
    .X(net656));
 clkbuf_2 fanout657 (.A(net658),
    .X(net657));
 dlymetal6s2s_1 fanout658 (.A(net662),
    .X(net658));
 clkbuf_2 fanout659 (.A(net660),
    .X(net659));
 clkbuf_2 fanout660 (.A(net662),
    .X(net660));
 clkbuf_2 fanout661 (.A(net662),
    .X(net661));
 clkbuf_2 fanout662 (.A(net675),
    .X(net662));
 clkbuf_2 fanout663 (.A(net665),
    .X(net663));
 clkbuf_2 fanout664 (.A(net667),
    .X(net664));
 dlymetal6s2s_1 fanout665 (.A(net667),
    .X(net665));
 clkbuf_2 fanout666 (.A(net667),
    .X(net666));
 clkbuf_2 fanout667 (.A(net675),
    .X(net667));
 clkbuf_2 fanout668 (.A(net669),
    .X(net668));
 dlymetal6s2s_1 fanout669 (.A(net675),
    .X(net669));
 clkbuf_2 fanout670 (.A(net675),
    .X(net670));
 clkbuf_2 fanout671 (.A(net674),
    .X(net671));
 clkbuf_2 fanout672 (.A(net674),
    .X(net672));
 clkbuf_1 fanout673 (.A(net674),
    .X(net673));
 clkbuf_2 fanout674 (.A(net675),
    .X(net674));
 buf_2 fanout675 (.A(_06407_),
    .X(net675));
 buf_2 fanout676 (.A(net677),
    .X(net676));
 buf_2 fanout677 (.A(_06303_),
    .X(net677));
 clkbuf_4 fanout678 (.A(net679),
    .X(net678));
 clkbuf_4 fanout679 (.A(_04419_),
    .X(net679));
 clkbuf_4 fanout680 (.A(net681),
    .X(net680));
 buf_2 fanout681 (.A(_02654_),
    .X(net681));
 buf_2 fanout682 (.A(_11403_),
    .X(net682));
 buf_2 fanout683 (.A(_11396_),
    .X(net683));
 buf_2 fanout684 (.A(net685),
    .X(net684));
 clkbuf_2 fanout685 (.A(net692),
    .X(net685));
 buf_2 fanout686 (.A(net688),
    .X(net686));
 buf_1 fanout687 (.A(net688),
    .X(net687));
 buf_2 fanout688 (.A(net692),
    .X(net688));
 buf_2 fanout689 (.A(net691),
    .X(net689));
 buf_2 fanout690 (.A(net691),
    .X(net690));
 clkbuf_2 fanout691 (.A(net692),
    .X(net691));
 clkbuf_2 fanout692 (.A(_07164_),
    .X(net692));
 buf_2 fanout693 (.A(net695),
    .X(net693));
 buf_2 fanout694 (.A(net695),
    .X(net694));
 clkbuf_2 fanout695 (.A(_07164_),
    .X(net695));
 buf_2 fanout696 (.A(net698),
    .X(net696));
 clkbuf_2 fanout697 (.A(_07164_),
    .X(net697));
 buf_2 fanout698 (.A(_07164_),
    .X(net698));
 buf_2 fanout699 (.A(net700),
    .X(net699));
 buf_2 fanout700 (.A(_07120_),
    .X(net700));
 clkbuf_2 fanout701 (.A(\digitop_pav2.sec_inst.shift_out.st[1] ),
    .X(net701));
 clkbuf_4 fanout702 (.A(\digitop_pav2.sec_inst.ld_mem.round_i ),
    .X(net702));
 clkbuf_2 fanout703 (.A(\digitop_pav2.sec_inst.shift_out.ctr[3] ),
    .X(net703));
 buf_1 fanout704 (.A(\digitop_pav2.sec_inst.shift_out.ctr[3] ),
    .X(net704));
 clkbuf_2 fanout705 (.A(net706),
    .X(net705));
 clkbuf_2 fanout706 (.A(\digitop_pav2.sec_inst.shift_out.ctr[2] ),
    .X(net706));
 clkbuf_2 fanout707 (.A(\digitop_pav2.sec_inst.shift_out.st[6] ),
    .X(net707));
 buf_2 fanout708 (.A(\digitop_pav2.sec_inst.shift_out.st[3] ),
    .X(net708));
 buf_2 fanout709 (.A(\digitop_pav2.sec_inst.shift_out.st[3] ),
    .X(net709));
 clkbuf_4 fanout710 (.A(net711),
    .X(net710));
 clkbuf_4 fanout711 (.A(\digitop_pav2.sec_inst.en_reg128 ),
    .X(net711));
 clkbuf_4 fanout712 (.A(net713),
    .X(net712));
 buf_2 fanout713 (.A(\digitop_pav2.sec_inst.en_reg128 ),
    .X(net713));
 buf_2 fanout714 (.A(\digitop_pav2.sec_inst.dg_key.en_i ),
    .X(net714));
 clkbuf_4 fanout715 (.A(\digitop_pav2.sec_inst.en_ld_data ),
    .X(net715));
 buf_2 fanout716 (.A(net717),
    .X(net716));
 clkbuf_2 fanout717 (.A(net718),
    .X(net717));
 clkbuf_2 fanout718 (.A(net719),
    .X(net718));
 dlymetal6s2s_1 fanout719 (.A(\digitop_pav2.sec_inst.en_ld_r ),
    .X(net719));
 clkbuf_2 fanout720 (.A(net722),
    .X(net720));
 clkbuf_2 fanout721 (.A(net722),
    .X(net721));
 clkbuf_2 fanout722 (.A(net723),
    .X(net722));
 buf_2 fanout723 (.A(net729),
    .X(net723));
 clkbuf_2 fanout724 (.A(net726),
    .X(net724));
 clkbuf_2 fanout725 (.A(net726),
    .X(net725));
 clkbuf_2 fanout726 (.A(net729),
    .X(net726));
 clkbuf_2 fanout727 (.A(net729),
    .X(net727));
 buf_1 fanout728 (.A(net729),
    .X(net728));
 clkbuf_2 fanout729 (.A(_03766_),
    .X(net729));
 clkbuf_2 fanout730 (.A(net732),
    .X(net730));
 clkbuf_2 fanout731 (.A(net732),
    .X(net731));
 dlymetal6s2s_1 fanout732 (.A(net757),
    .X(net732));
 clkbuf_2 fanout733 (.A(net757),
    .X(net733));
 clkbuf_2 fanout734 (.A(net757),
    .X(net734));
 clkbuf_2 fanout735 (.A(net742),
    .X(net735));
 buf_1 fanout736 (.A(net742),
    .X(net736));
 clkbuf_2 fanout737 (.A(net742),
    .X(net737));
 clkbuf_2 fanout738 (.A(net742),
    .X(net738));
 clkbuf_2 fanout739 (.A(net742),
    .X(net739));
 clkbuf_2 fanout740 (.A(net742),
    .X(net740));
 buf_1 fanout741 (.A(net742),
    .X(net741));
 clkbuf_4 fanout742 (.A(net757),
    .X(net742));
 clkbuf_2 fanout743 (.A(net745),
    .X(net743));
 clkbuf_2 fanout744 (.A(net745),
    .X(net744));
 clkbuf_2 fanout745 (.A(net757),
    .X(net745));
 clkbuf_2 fanout746 (.A(net748),
    .X(net746));
 buf_1 fanout747 (.A(net748),
    .X(net747));
 buf_1 fanout748 (.A(net757),
    .X(net748));
 clkbuf_2 fanout749 (.A(net752),
    .X(net749));
 clkbuf_2 fanout750 (.A(net752),
    .X(net750));
 buf_1 fanout751 (.A(net752),
    .X(net751));
 dlymetal6s2s_1 fanout752 (.A(net757),
    .X(net752));
 clkbuf_2 fanout753 (.A(net756),
    .X(net753));
 clkbuf_2 fanout754 (.A(net755),
    .X(net754));
 clkbuf_2 fanout755 (.A(net756),
    .X(net755));
 clkbuf_2 fanout756 (.A(net757),
    .X(net756));
 clkbuf_4 fanout757 (.A(_03766_),
    .X(net757));
 clkbuf_2 fanout758 (.A(net759),
    .X(net758));
 clkbuf_2 fanout759 (.A(net761),
    .X(net759));
 buf_2 fanout760 (.A(net761),
    .X(net760));
 dlymetal6s2s_1 fanout761 (.A(net762),
    .X(net761));
 buf_2 fanout762 (.A(net769),
    .X(net762));
 clkbuf_2 fanout763 (.A(net765),
    .X(net763));
 clkbuf_2 fanout764 (.A(net765),
    .X(net764));
 buf_2 fanout765 (.A(net768),
    .X(net765));
 clkbuf_2 fanout766 (.A(net768),
    .X(net766));
 clkbuf_2 fanout767 (.A(net768),
    .X(net767));
 clkbuf_2 fanout768 (.A(net769),
    .X(net768));
 buf_2 fanout769 (.A(_03765_),
    .X(net769));
 clkbuf_2 fanout770 (.A(net776),
    .X(net770));
 buf_1 fanout771 (.A(net776),
    .X(net771));
 buf_2 fanout772 (.A(net776),
    .X(net772));
 buf_1 fanout773 (.A(net776),
    .X(net773));
 buf_2 fanout774 (.A(net775),
    .X(net774));
 clkbuf_2 fanout775 (.A(net776),
    .X(net775));
 clkbuf_2 fanout776 (.A(net800),
    .X(net776));
 clkbuf_2 fanout777 (.A(net785),
    .X(net777));
 dlymetal6s2s_1 fanout778 (.A(net785),
    .X(net778));
 clkbuf_2 fanout779 (.A(net785),
    .X(net779));
 clkbuf_1 fanout780 (.A(net785),
    .X(net780));
 buf_2 fanout781 (.A(net784),
    .X(net781));
 clkbuf_2 fanout782 (.A(net783),
    .X(net782));
 clkbuf_2 fanout783 (.A(net784),
    .X(net783));
 clkbuf_2 fanout784 (.A(net785),
    .X(net784));
 clkbuf_2 fanout785 (.A(net800),
    .X(net785));
 buf_2 fanout786 (.A(net788),
    .X(net786));
 clkbuf_2 fanout787 (.A(net788),
    .X(net787));
 clkbuf_2 fanout788 (.A(net800),
    .X(net788));
 clkbuf_2 fanout789 (.A(net791),
    .X(net789));
 buf_1 fanout790 (.A(net791),
    .X(net790));
 dlymetal6s2s_1 fanout791 (.A(net800),
    .X(net791));
 buf_2 fanout792 (.A(net795),
    .X(net792));
 clkbuf_2 fanout793 (.A(net795),
    .X(net793));
 clkbuf_2 fanout794 (.A(net795),
    .X(net794));
 clkbuf_2 fanout795 (.A(net800),
    .X(net795));
 clkbuf_2 fanout796 (.A(net799),
    .X(net796));
 clkbuf_2 fanout797 (.A(net799),
    .X(net797));
 buf_1 fanout798 (.A(net799),
    .X(net798));
 clkbuf_2 fanout799 (.A(net800),
    .X(net799));
 clkbuf_4 fanout800 (.A(net801),
    .X(net800));
 buf_1 wire801 (.A(_03765_),
    .X(net801));
 clkbuf_2 wire802 (.A(_03661_),
    .X(net802));
 buf_2 fanout803 (.A(_08107_),
    .X(net803));
 buf_2 fanout804 (.A(net805),
    .X(net804));
 buf_2 fanout805 (.A(_08106_),
    .X(net805));
 clkbuf_4 fanout806 (.A(net807),
    .X(net806));
 buf_2 fanout807 (.A(_07450_),
    .X(net807));
 buf_2 fanout808 (.A(_07337_),
    .X(net808));
 buf_2 fanout809 (.A(_05262_),
    .X(net809));
 buf_2 fanout810 (.A(_05262_),
    .X(net810));
 clkbuf_4 fanout811 (.A(_07603_),
    .X(net811));
 buf_2 fanout812 (.A(net1641),
    .X(net812));
 clkbuf_2 fanout813 (.A(net1640),
    .X(net813));
 clkbuf_2 fanout814 (.A(net815),
    .X(net814));
 clkbuf_2 fanout815 (.A(net816),
    .X(net815));
 clkbuf_2 fanout816 (.A(net1640),
    .X(net816));
 clkbuf_4 fanout817 (.A(net1639),
    .X(net817));
 clkbuf_4 fanout818 (.A(net819),
    .X(net818));
 buf_4 fanout819 (.A(net1645),
    .X(net819));
 clkbuf_2 fanout820 (.A(net821),
    .X(net820));
 clkbuf_2 fanout821 (.A(net822),
    .X(net821));
 clkbuf_2 fanout822 (.A(net823),
    .X(net822));
 clkbuf_2 fanout823 (.A(net829),
    .X(net823));
 clkbuf_2 fanout824 (.A(net825),
    .X(net824));
 buf_1 fanout825 (.A(net826),
    .X(net825));
 clkbuf_2 fanout826 (.A(net828),
    .X(net826));
 clkbuf_2 fanout827 (.A(net828),
    .X(net827));
 clkbuf_2 fanout828 (.A(net829),
    .X(net828));
 buf_2 fanout829 (.A(_06763_),
    .X(net829));
 clkbuf_2 fanout830 (.A(net831),
    .X(net830));
 clkbuf_2 fanout831 (.A(net832),
    .X(net831));
 clkbuf_2 fanout832 (.A(net841),
    .X(net832));
 clkbuf_2 fanout833 (.A(net841),
    .X(net833));
 buf_1 fanout834 (.A(net841),
    .X(net834));
 clkbuf_2 fanout835 (.A(net837),
    .X(net835));
 clkbuf_2 fanout836 (.A(net841),
    .X(net836));
 buf_1 fanout837 (.A(net841),
    .X(net837));
 clkbuf_2 fanout838 (.A(net840),
    .X(net838));
 clkbuf_2 fanout839 (.A(net840),
    .X(net839));
 clkbuf_2 fanout840 (.A(net841),
    .X(net840));
 buf_2 fanout841 (.A(_06763_),
    .X(net841));
 clkbuf_2 fanout842 (.A(net843),
    .X(net842));
 buf_2 fanout843 (.A(net852),
    .X(net843));
 clkbuf_2 fanout844 (.A(net845),
    .X(net844));
 clkbuf_2 fanout845 (.A(net852),
    .X(net845));
 clkbuf_2 fanout846 (.A(net851),
    .X(net846));
 clkbuf_2 fanout847 (.A(net848),
    .X(net847));
 clkbuf_2 fanout848 (.A(net851),
    .X(net848));
 clkbuf_2 fanout849 (.A(net850),
    .X(net849));
 clkbuf_2 fanout850 (.A(net851),
    .X(net850));
 buf_2 fanout851 (.A(net852),
    .X(net851));
 clkbuf_2 fanout852 (.A(_06763_),
    .X(net852));
 clkbuf_2 fanout853 (.A(net855),
    .X(net853));
 clkbuf_2 fanout854 (.A(net855),
    .X(net854));
 clkbuf_2 fanout855 (.A(net856),
    .X(net855));
 clkbuf_2 fanout856 (.A(_06411_),
    .X(net856));
 clkbuf_2 fanout857 (.A(net858),
    .X(net857));
 buf_2 fanout858 (.A(net861),
    .X(net858));
 clkbuf_2 fanout859 (.A(net861),
    .X(net859));
 buf_1 fanout860 (.A(net861),
    .X(net860));
 clkbuf_2 fanout861 (.A(_06411_),
    .X(net861));
 clkbuf_2 fanout862 (.A(net886),
    .X(net862));
 buf_1 fanout863 (.A(net886),
    .X(net863));
 clkbuf_2 fanout864 (.A(net865),
    .X(net864));
 clkbuf_2 fanout865 (.A(net886),
    .X(net865));
 clkbuf_2 fanout866 (.A(net873),
    .X(net866));
 dlymetal6s2s_1 fanout867 (.A(net873),
    .X(net867));
 clkbuf_2 fanout868 (.A(net873),
    .X(net868));
 buf_1 fanout869 (.A(net873),
    .X(net869));
 clkbuf_2 fanout870 (.A(net872),
    .X(net870));
 buf_1 fanout871 (.A(net872),
    .X(net871));
 buf_2 fanout872 (.A(net873),
    .X(net872));
 clkbuf_2 fanout873 (.A(net886),
    .X(net873));
 clkbuf_2 fanout874 (.A(net876),
    .X(net874));
 clkbuf_2 fanout875 (.A(net876),
    .X(net875));
 clkbuf_2 fanout876 (.A(net886),
    .X(net876));
 clkbuf_2 fanout877 (.A(net878),
    .X(net877));
 buf_1 fanout878 (.A(net886),
    .X(net878));
 clkbuf_2 fanout879 (.A(net885),
    .X(net879));
 clkbuf_2 fanout880 (.A(net885),
    .X(net880));
 clkbuf_2 fanout881 (.A(net882),
    .X(net881));
 clkbuf_2 fanout882 (.A(net884),
    .X(net882));
 clkbuf_2 fanout883 (.A(net884),
    .X(net883));
 dlymetal6s2s_1 fanout884 (.A(net885),
    .X(net884));
 clkbuf_2 fanout885 (.A(net886),
    .X(net885));
 clkbuf_4 fanout886 (.A(_06411_),
    .X(net886));
 clkbuf_4 fanout887 (.A(net889),
    .X(net887));
 clkbuf_2 fanout888 (.A(net889),
    .X(net888));
 buf_2 fanout889 (.A(net892),
    .X(net889));
 clkbuf_4 fanout890 (.A(net891),
    .X(net890));
 buf_4 fanout891 (.A(net892),
    .X(net891));
 buf_2 fanout892 (.A(_03760_),
    .X(net892));
 clkbuf_4 fanout893 (.A(net895),
    .X(net893));
 clkbuf_2 fanout894 (.A(net895),
    .X(net894));
 clkbuf_4 fanout895 (.A(net905),
    .X(net895));
 clkbuf_4 fanout896 (.A(net899),
    .X(net896));
 clkbuf_4 fanout897 (.A(net899),
    .X(net897));
 clkbuf_2 fanout898 (.A(net899),
    .X(net898));
 buf_2 fanout899 (.A(net905),
    .X(net899));
 clkbuf_4 fanout900 (.A(net901),
    .X(net900));
 buf_4 fanout901 (.A(net905),
    .X(net901));
 clkbuf_4 fanout902 (.A(net904),
    .X(net902));
 clkbuf_4 fanout903 (.A(net904),
    .X(net903));
 clkbuf_4 fanout904 (.A(net905),
    .X(net904));
 clkbuf_4 fanout905 (.A(_03760_),
    .X(net905));
 buf_4 fanout906 (.A(_03759_),
    .X(net906));
 clkbuf_4 fanout907 (.A(net908),
    .X(net907));
 clkbuf_4 fanout908 (.A(net911),
    .X(net908));
 buf_2 fanout909 (.A(net910),
    .X(net909));
 buf_4 fanout910 (.A(net911),
    .X(net910));
 clkbuf_4 fanout911 (.A(_03759_),
    .X(net911));
 clkbuf_4 fanout912 (.A(_07528_),
    .X(net912));
 clkbuf_4 fanout913 (.A(_07527_),
    .X(net913));
 clkbuf_4 fanout914 (.A(_04907_),
    .X(net914));
 buf_2 fanout915 (.A(_04907_),
    .X(net915));
 clkbuf_4 fanout916 (.A(net918),
    .X(net916));
 clkbuf_4 fanout917 (.A(net918),
    .X(net917));
 clkbuf_4 fanout918 (.A(net919),
    .X(net918));
 clkbuf_4 fanout919 (.A(net924),
    .X(net919));
 clkbuf_4 fanout920 (.A(net922),
    .X(net920));
 clkbuf_4 fanout921 (.A(net922),
    .X(net921));
 clkbuf_2 fanout922 (.A(net923),
    .X(net922));
 buf_2 fanout923 (.A(net924),
    .X(net923));
 buf_2 fanout924 (.A(_03762_),
    .X(net924));
 clkbuf_4 fanout925 (.A(net930),
    .X(net925));
 clkbuf_2 fanout926 (.A(net930),
    .X(net926));
 clkbuf_4 fanout927 (.A(net930),
    .X(net927));
 clkbuf_4 fanout928 (.A(net929),
    .X(net928));
 clkbuf_4 fanout929 (.A(net930),
    .X(net929));
 clkbuf_2 fanout930 (.A(net951),
    .X(net930));
 clkbuf_4 fanout931 (.A(net938),
    .X(net931));
 clkbuf_4 fanout932 (.A(net938),
    .X(net932));
 clkbuf_2 fanout933 (.A(net938),
    .X(net933));
 clkbuf_4 fanout934 (.A(net937),
    .X(net934));
 clkbuf_4 fanout935 (.A(net937),
    .X(net935));
 clkbuf_2 fanout936 (.A(net937),
    .X(net936));
 clkbuf_2 fanout937 (.A(net938),
    .X(net937));
 clkbuf_2 fanout938 (.A(net951),
    .X(net938));
 clkbuf_4 fanout939 (.A(net941),
    .X(net939));
 clkbuf_4 fanout940 (.A(net941),
    .X(net940));
 clkbuf_2 fanout941 (.A(net951),
    .X(net941));
 clkbuf_4 fanout942 (.A(net943),
    .X(net942));
 clkbuf_4 fanout943 (.A(net951),
    .X(net943));
 clkbuf_4 fanout944 (.A(net946),
    .X(net944));
 clkbuf_4 fanout945 (.A(net946),
    .X(net945));
 buf_2 fanout946 (.A(net951),
    .X(net946));
 clkbuf_4 fanout947 (.A(net950),
    .X(net947));
 clkbuf_4 fanout948 (.A(net950),
    .X(net948));
 clkbuf_2 fanout949 (.A(net950),
    .X(net949));
 clkbuf_2 fanout950 (.A(net951),
    .X(net950));
 clkbuf_4 fanout951 (.A(_03762_),
    .X(net951));
 clkbuf_4 fanout952 (.A(net955),
    .X(net952));
 buf_4 fanout953 (.A(net955),
    .X(net953));
 buf_2 fanout954 (.A(net955),
    .X(net954));
 clkbuf_4 fanout955 (.A(_03761_),
    .X(net955));
 buf_2 fanout956 (.A(_09416_),
    .X(net956));
 buf_2 fanout957 (.A(_09389_),
    .X(net957));
 buf_2 fanout958 (.A(_08113_),
    .X(net958));
 buf_2 fanout959 (.A(_08112_),
    .X(net959));
 buf_2 fanout960 (.A(net961),
    .X(net960));
 clkbuf_2 fanout961 (.A(_08110_),
    .X(net961));
 clkbuf_4 fanout962 (.A(_07508_),
    .X(net962));
 buf_4 fanout963 (.A(_07488_),
    .X(net963));
 clkbuf_4 fanout964 (.A(net965),
    .X(net964));
 clkbuf_4 fanout965 (.A(_07487_),
    .X(net965));
 buf_1 max_cap966 (.A(_07487_),
    .X(net966));
 buf_2 fanout967 (.A(net968),
    .X(net967));
 buf_2 fanout968 (.A(_07162_),
    .X(net968));
 buf_2 fanout969 (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.pro_abort_b_i ),
    .X(net969));
 clkbuf_4 fanout970 (.A(net971),
    .X(net970));
 buf_2 fanout971 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.ebv_en ),
    .X(net971));
 clkbuf_4 fanout972 (.A(net973),
    .X(net972));
 buf_2 fanout973 (.A(net1809),
    .X(net973));
 clkbuf_2 fanout974 (.A(_08965_),
    .X(net974));
 dlymetal6s2s_1 fanout975 (.A(_08965_),
    .X(net975));
 buf_2 fanout976 (.A(_08132_),
    .X(net976));
 clkbuf_2 fanout977 (.A(_08132_),
    .X(net977));
 buf_2 fanout978 (.A(net979),
    .X(net978));
 buf_2 fanout979 (.A(_08130_),
    .X(net979));
 clkbuf_4 fanout980 (.A(net981),
    .X(net980));
 clkbuf_2 fanout981 (.A(net983),
    .X(net981));
 clkbuf_4 fanout982 (.A(net983),
    .X(net982));
 clkbuf_2 fanout983 (.A(net1620),
    .X(net983));
 clkbuf_4 fanout984 (.A(net986),
    .X(net984));
 clkbuf_4 fanout985 (.A(net986),
    .X(net985));
 buf_2 fanout986 (.A(net1620),
    .X(net986));
 clkbuf_4 fanout987 (.A(net990),
    .X(net987));
 clkbuf_4 fanout988 (.A(net990),
    .X(net988));
 buf_2 fanout989 (.A(net990),
    .X(net989));
 dlymetal6s2s_1 fanout990 (.A(net1001),
    .X(net990));
 clkbuf_4 fanout991 (.A(net1001),
    .X(net991));
 buf_2 fanout992 (.A(net1001),
    .X(net992));
 clkbuf_4 fanout993 (.A(net996),
    .X(net993));
 clkbuf_4 fanout994 (.A(net996),
    .X(net994));
 clkbuf_2 fanout995 (.A(net996),
    .X(net995));
 dlymetal6s2s_1 fanout996 (.A(net1001),
    .X(net996));
 clkbuf_4 fanout997 (.A(net1000),
    .X(net997));
 clkbuf_4 fanout998 (.A(net1000),
    .X(net998));
 clkbuf_2 fanout999 (.A(net1000),
    .X(net999));
 clkbuf_2 fanout1000 (.A(net1001),
    .X(net1000));
 clkbuf_2 fanout1001 (.A(net1620),
    .X(net1001));
 clkbuf_4 fanout1002 (.A(net1003),
    .X(net1002));
 clkbuf_4 fanout1003 (.A(net1004),
    .X(net1003));
 clkbuf_4 fanout1004 (.A(net1620),
    .X(net1004));
 clkbuf_4 fanout1005 (.A(net1621),
    .X(net1005));
 clkbuf_2 fanout1006 (.A(net1621),
    .X(net1006));
 clkbuf_2 fanout1007 (.A(net1620),
    .X(net1007));
 clkbuf_4 fanout1008 (.A(net1619),
    .X(net1008));
 buf_2 fanout1009 (.A(net1010),
    .X(net1009));
 clkbuf_2 fanout1010 (.A(_07408_),
    .X(net1010));
 buf_2 fanout1011 (.A(_07343_),
    .X(net1011));
 buf_2 fanout1012 (.A(_03684_),
    .X(net1012));
 dlymetal6s2s_1 fanout1013 (.A(_03684_),
    .X(net1013));
 buf_2 fanout1014 (.A(_10325_),
    .X(net1014));
 buf_1 wire1015 (.A(_09022_),
    .X(net1015));
 buf_2 fanout1016 (.A(_07962_),
    .X(net1016));
 clkbuf_4 fanout1017 (.A(_07492_),
    .X(net1017));
 buf_1 wire1018 (.A(_07341_),
    .X(net1018));
 buf_2 fanout1019 (.A(_06153_),
    .X(net1019));
 buf_2 fanout1020 (.A(net1021),
    .X(net1020));
 buf_2 fanout1021 (.A(_04911_),
    .X(net1021));
 clkbuf_4 fanout1022 (.A(_04743_),
    .X(net1022));
 clkbuf_2 fanout1023 (.A(_10818_),
    .X(net1023));
 clkbuf_2 fanout1024 (.A(_10814_),
    .X(net1024));
 clkbuf_2 fanout1025 (.A(_09397_),
    .X(net1025));
 clkbuf_4 fanout1026 (.A(net1027),
    .X(net1026));
 clkbuf_2 fanout1027 (.A(_09385_),
    .X(net1027));
 clkbuf_4 fanout1028 (.A(_08046_),
    .X(net1028));
 buf_2 fanout1029 (.A(_08046_),
    .X(net1029));
 buf_4 max_cap1030 (.A(_07898_),
    .X(net1030));
 buf_2 fanout1031 (.A(_07617_),
    .X(net1031));
 buf_2 fanout1032 (.A(_07617_),
    .X(net1032));
 buf_4 fanout1033 (.A(_07577_),
    .X(net1033));
 clkbuf_2 max_cap1034 (.A(_07482_),
    .X(net1034));
 clkbuf_8 fanout1035 (.A(_07081_),
    .X(net1035));
 clkbuf_4 fanout1036 (.A(_07050_),
    .X(net1036));
 clkbuf_4 fanout1037 (.A(_07039_),
    .X(net1037));
 buf_2 fanout1038 (.A(_07035_),
    .X(net1038));
 clkbuf_2 fanout1039 (.A(_07035_),
    .X(net1039));
 clkbuf_2 fanout1040 (.A(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[3] ),
    .X(net1040));
 clkbuf_2 fanout1041 (.A(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[3] ),
    .X(net1041));
 buf_2 fanout1042 (.A(\digitop_pav2.access_inst.access_transceiver0.dt_ptr[2] ),
    .X(net1042));
 clkbuf_4 fanout1043 (.A(net1044),
    .X(net1043));
 clkbuf_2 fanout1044 (.A(net1045),
    .X(net1044));
 buf_2 fanout1045 (.A(\digitop_pav2.access_inst.access_transceiver0.ctrl_circ_buf ),
    .X(net1045));
 buf_2 fanout1046 (.A(net1048),
    .X(net1046));
 buf_1 fanout1047 (.A(net1048),
    .X(net1047));
 clkbuf_4 fanout1048 (.A(\digitop_pav2.access_inst.access_ctrl0.proc_finish0_i ),
    .X(net1048));
 buf_2 fanout1049 (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[0] ),
    .X(net1049));
 clkbuf_2 fanout1050 (.A(net1051),
    .X(net1050));
 buf_2 fanout1051 (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[8] ),
    .X(net1051));
 clkbuf_2 fanout1052 (.A(net1053),
    .X(net1052));
 buf_2 fanout1053 (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[7] ),
    .X(net1053));
 buf_2 fanout1054 (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[3] ),
    .X(net1054));
 buf_1 fanout1055 (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[3] ),
    .X(net1055));
 clkbuf_4 fanout1056 (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[2] ),
    .X(net1056));
 buf_1 fanout1057 (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[2] ),
    .X(net1057));
 buf_2 fanout1058 (.A(net1059),
    .X(net1058));
 clkbuf_2 fanout1059 (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[1] ),
    .X(net1059));
 buf_2 fanout1060 (.A(net1061),
    .X(net1060));
 clkbuf_2 fanout1061 (.A(net1062),
    .X(net1061));
 clkbuf_2 fanout1062 (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[0] ),
    .X(net1062));
 clkbuf_4 fanout1063 (.A(\digitop_pav2.access_inst.access_ctrl0.ld_dt_env_finish_i ),
    .X(net1063));
 clkbuf_2 fanout1064 (.A(\digitop_pav2.access_inst.access_ctrl0.ld_dt_env_finish_i ),
    .X(net1064));
 buf_2 fanout1065 (.A(\digitop_pav2.access_inst.access_check0.proc_finish1_i ),
    .X(net1065));
 buf_2 fanout1066 (.A(\digitop_pav2.access_inst.access_ctrl0.wr_key_finish_i ),
    .X(net1066));
 buf_1 fanout1067 (.A(\digitop_pav2.access_inst.access_ctrl0.wr_key_finish_i ),
    .X(net1067));
 buf_2 fanout1068 (.A(net1070),
    .X(net1068));
 buf_2 fanout1069 (.A(net1070),
    .X(net1069));
 clkbuf_2 fanout1070 (.A(\digitop_pav2.access_inst.access_check0.wr_check_sync_o ),
    .X(net1070));
 clkbuf_4 fanout1071 (.A(\digitop_pav2.access_inst.access_check0.wcnt_check_one ),
    .X(net1071));
 clkbuf_4 fanout1072 (.A(\digitop_pav2.access_inst.access_check0.wordptr_i[6] ),
    .X(net1072));
 buf_2 fanout1073 (.A(\digitop_pav2.access_inst.access_check0.wordptr_i[5] ),
    .X(net1073));
 buf_2 fanout1074 (.A(\digitop_pav2.access_inst.access_check0.wordptr_i[4] ),
    .X(net1074));
 clkbuf_2 fanout1075 (.A(net1076),
    .X(net1075));
 buf_2 fanout1076 (.A(\digitop_pav2.access_inst.access_check0.wordptr_i[3] ),
    .X(net1076));
 clkbuf_2 fanout1077 (.A(net1078),
    .X(net1077));
 buf_2 fanout1078 (.A(\digitop_pav2.access_inst.access_check0.wordptr_i[2] ),
    .X(net1078));
 clkbuf_2 fanout1079 (.A(net1080),
    .X(net1079));
 buf_2 fanout1080 (.A(\digitop_pav2.access_inst.access_check0.wordptr_i[1] ),
    .X(net1080));
 buf_2 fanout1081 (.A(net1082),
    .X(net1081));
 dlymetal6s2s_1 fanout1082 (.A(\digitop_pav2.access_inst.access_check0.wordptr_i[0] ),
    .X(net1082));
 clkbuf_4 fanout1083 (.A(net1085),
    .X(net1083));
 buf_2 fanout1084 (.A(net1085),
    .X(net1084));
 buf_2 fanout1085 (.A(net1086),
    .X(net1085));
 buf_4 fanout1086 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[15] ),
    .X(net1086));
 buf_4 fanout1087 (.A(net1088),
    .X(net1087));
 buf_2 fanout1088 (.A(net1089),
    .X(net1088));
 clkbuf_4 fanout1089 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[14] ),
    .X(net1089));
 clkbuf_4 fanout1090 (.A(net1092),
    .X(net1090));
 buf_2 fanout1091 (.A(net1092),
    .X(net1091));
 buf_2 fanout1092 (.A(net1093),
    .X(net1092));
 buf_4 fanout1093 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[13] ),
    .X(net1093));
 buf_4 fanout1094 (.A(net1095),
    .X(net1094));
 buf_4 fanout1095 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[12] ),
    .X(net1095));
 buf_4 fanout1096 (.A(net1097),
    .X(net1096));
 buf_4 fanout1097 (.A(net1098),
    .X(net1097));
 buf_4 fanout1098 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[11] ),
    .X(net1098));
 buf_4 fanout1099 (.A(net1101),
    .X(net1099));
 clkbuf_2 fanout1100 (.A(net1101),
    .X(net1100));
 clkbuf_4 fanout1101 (.A(net1102),
    .X(net1101));
 buf_4 fanout1102 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[10] ),
    .X(net1102));
 clkbuf_4 fanout1103 (.A(net1105),
    .X(net1103));
 buf_2 fanout1104 (.A(net1105),
    .X(net1104));
 clkbuf_4 fanout1105 (.A(net1106),
    .X(net1105));
 clkbuf_8 fanout1106 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[9] ),
    .X(net1106));
 buf_4 fanout1107 (.A(net1109),
    .X(net1107));
 clkbuf_2 fanout1108 (.A(net1109),
    .X(net1108));
 buf_2 fanout1109 (.A(net1110),
    .X(net1109));
 clkbuf_4 fanout1110 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[8] ),
    .X(net1110));
 clkbuf_4 fanout1111 (.A(net1112),
    .X(net1111));
 buf_2 fanout1112 (.A(net1113),
    .X(net1112));
 clkbuf_4 fanout1113 (.A(net1114),
    .X(net1113));
 clkbuf_8 fanout1114 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[7] ),
    .X(net1114));
 buf_4 fanout1115 (.A(net1116),
    .X(net1115));
 buf_2 fanout1116 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[6] ),
    .X(net1116));
 buf_4 fanout1117 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[6] ),
    .X(net1117));
 buf_4 fanout1118 (.A(net1119),
    .X(net1118));
 clkbuf_4 fanout1119 (.A(net1120),
    .X(net1119));
 clkbuf_4 fanout1120 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[5] ),
    .X(net1120));
 buf_4 fanout1121 (.A(net1122),
    .X(net1121));
 buf_2 fanout1122 (.A(net1123),
    .X(net1122));
 buf_4 fanout1123 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[4] ),
    .X(net1123));
 clkbuf_4 fanout1124 (.A(net1125),
    .X(net1124));
 buf_2 fanout1125 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[3] ),
    .X(net1125));
 buf_4 fanout1126 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[3] ),
    .X(net1126));
 buf_4 fanout1127 (.A(net1129),
    .X(net1127));
 clkbuf_2 fanout1128 (.A(net1129),
    .X(net1128));
 buf_2 fanout1129 (.A(net1130),
    .X(net1129));
 clkbuf_4 fanout1130 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[2] ),
    .X(net1130));
 buf_4 fanout1131 (.A(net1133),
    .X(net1131));
 buf_4 fanout1132 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[1] ),
    .X(net1132));
 clkbuf_4 fanout1133 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[1] ),
    .X(net1133));
 buf_4 fanout1134 (.A(net1135),
    .X(net1134));
 buf_6 fanout1135 (.A(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[0] ),
    .X(net1135));
 buf_2 fanout1136 (.A(net1137),
    .X(net1136));
 buf_2 fanout1137 (.A(net1138),
    .X(net1137));
 buf_2 fanout1138 (.A(\digitop_pav2.memctrl_inst.addr_to_reram[4] ),
    .X(net1138));
 buf_2 fanout1139 (.A(net1141),
    .X(net1139));
 buf_2 fanout1140 (.A(net1141),
    .X(net1140));
 buf_2 fanout1141 (.A(\digitop_pav2.memctrl_inst.addr_to_reram[3] ),
    .X(net1141));
 buf_2 fanout1142 (.A(\digitop_pav2.access_inst.access_ctrl0.state[25] ),
    .X(net1142));
 buf_2 fanout1143 (.A(\digitop_pav2.access_inst.access_ctrl0.state[19] ),
    .X(net1143));
 clkbuf_4 fanout1144 (.A(\digitop_pav2.access_inst.access_ctrl0.ctrl_ld_dt_ok ),
    .X(net1144));
 clkbuf_4 fanout1145 (.A(\digitop_pav2.access_inst.access_ctrl0.crc_en_o ),
    .X(net1145));
 buf_2 fanout1146 (.A(net1147),
    .X(net1146));
 buf_2 fanout1147 (.A(net1148),
    .X(net1147));
 buf_2 fanout1148 (.A(\digitop_pav2.access_inst.access_check0.wr_key_ck_i ),
    .X(net1148));
 buf_2 fanout1149 (.A(\digitop_pav2.access_inst.access_check0.wr_key_ck_i ),
    .X(net1149));
 clkbuf_2 fanout1150 (.A(\digitop_pav2.access_inst.access_check0.wr_key_ck_i ),
    .X(net1150));
 buf_2 fanout1151 (.A(\digitop_pav2.access_inst.access_check0.write_check_i ),
    .X(net1151));
 dlymetal6s2s_1 fanout1152 (.A(\digitop_pav2.access_inst.access_check0.write_check_i ),
    .X(net1152));
 clkbuf_4 fanout1153 (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[2] ),
    .X(net1153));
 clkbuf_2 fanout1154 (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[2] ),
    .X(net1154));
 clkbuf_4 fanout1155 (.A(\digitop_pav2.access_inst.access_proc0.proc_crc_check[2] ),
    .X(net1155));
 buf_2 fanout1156 (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[5] ),
    .X(net1156));
 buf_2 fanout1157 (.A(net1158),
    .X(net1157));
 buf_2 fanout1158 (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[4] ),
    .X(net1158));
 buf_2 fanout1159 (.A(\digitop_pav2.access_inst.access_proc0.nvm_acc_addr[6] ),
    .X(net1159));
 clkbuf_4 fanout1160 (.A(net1161),
    .X(net1160));
 buf_2 fanout1161 (.A(_06144_),
    .X(net1161));
 clkbuf_2 max_cap1162 (.A(_10461_),
    .X(net1162));
 clkbuf_2 max_cap1163 (.A(_09150_),
    .X(net1163));
 buf_2 fanout1164 (.A(net1165),
    .X(net1164));
 clkbuf_2 fanout1165 (.A(_07338_),
    .X(net1165));
 clkbuf_4 fanout1166 (.A(net1167),
    .X(net1166));
 buf_2 fanout1167 (.A(_07272_),
    .X(net1167));
 clkbuf_4 fanout1168 (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[2] ),
    .X(net1168));
 buf_2 fanout1169 (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.q[1] ),
    .X(net1169));
 buf_2 fanout1170 (.A(net1172),
    .X(net1170));
 dlymetal6s2s_1 fanout1171 (.A(net1172),
    .X(net1171));
 clkbuf_2 fanout1172 (.A(\digitop_pav2.invent_inst.invent_qqqr_pav2.state[2] ),
    .X(net1172));
 clkbuf_2 fanout1173 (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[3] ),
    .X(net1173));
 clkbuf_2 fanout1174 (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[2] ),
    .X(net1174));
 clkbuf_2 fanout1175 (.A(\digitop_pav2.invent_inst.invent_sel_pav2.bitptr[1] ),
    .X(net1175));
 clkbuf_2 fanout1176 (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[2] ),
    .X(net1176));
 clkbuf_2 fanout1177 (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_ctr_o[1] ),
    .X(net1177));
 clkbuf_4 fanout1178 (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer2_o[0] ),
    .X(net1178));
 buf_2 fanout1179 (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[2] ),
    .X(net1179));
 clkbuf_2 fanout1180 (.A(\digitop_pav2.invent_inst.invent_buffer_pav2.rx_buffer1_o[1] ),
    .X(net1180));
 buf_2 fanout1181 (.A(_07258_),
    .X(net1181));
 clkbuf_2 fanout1182 (.A(\digitop_pav2.ack_inst.cnt_ff[1] ),
    .X(net1182));
 clkbuf_2 max_cap1183 (.A(net1184),
    .X(net1183));
 clkbuf_2 wire1184 (.A(_07324_),
    .X(net1184));
 buf_2 fanout1185 (.A(_07305_),
    .X(net1185));
 clkbuf_4 fanout1186 (.A(_07243_),
    .X(net1186));
 clkbuf_2 max_cap1187 (.A(_09030_),
    .X(net1187));
 buf_2 fanout1188 (.A(_09016_),
    .X(net1188));
 clkbuf_2 fanout1189 (.A(_09016_),
    .X(net1189));
 clkbuf_4 fanout1190 (.A(net1193),
    .X(net1190));
 buf_2 fanout1191 (.A(net1193),
    .X(net1191));
 buf_1 fanout1192 (.A(net1193),
    .X(net1192));
 clkbuf_2 fanout1193 (.A(\digitop_pav2.sync_inst.inst_clkx.g_access ),
    .X(net1193));
 buf_2 fanout1194 (.A(\digitop_pav2.sync_inst.inst_clkx.g_access ),
    .X(net1194));
 clkbuf_4 fanout1195 (.A(_07310_),
    .X(net1195));
 buf_2 fanout1196 (.A(_07289_),
    .X(net1196));
 buf_2 fanout1197 (.A(_07269_),
    .X(net1197));
 buf_2 wire1198 (.A(_07247_),
    .X(net1198));
 buf_4 fanout1199 (.A(net1692),
    .X(net1199));
 buf_2 fanout1200 (.A(net1203),
    .X(net1200));
 buf_4 fanout1201 (.A(net1203),
    .X(net1201));
 buf_4 fanout1202 (.A(net1203),
    .X(net1202));
 buf_2 fanout1203 (.A(net1697),
    .X(net1203));
 clkbuf_4 fanout1204 (.A(net1205),
    .X(net1204));
 clkbuf_4 fanout1205 (.A(net1208),
    .X(net1205));
 clkbuf_4 fanout1206 (.A(net1208),
    .X(net1206));
 buf_2 fanout1207 (.A(net1208),
    .X(net1207));
 buf_2 fanout1208 (.A(net1212),
    .X(net1208));
 buf_4 fanout1209 (.A(net1212),
    .X(net1209));
 clkbuf_4 fanout1210 (.A(net1212),
    .X(net1210));
 clkbuf_2 fanout1211 (.A(net1212),
    .X(net1211));
 clkbuf_2 fanout1212 (.A(net1213),
    .X(net1212));
 buf_4 fanout1213 (.A(net1697),
    .X(net1213));
 buf_2 fanout1214 (.A(net1696),
    .X(net1214));
 clkbuf_4 fanout1215 (.A(net1216),
    .X(net1215));
 clkbuf_2 fanout1216 (.A(_07282_),
    .X(net1216));
 buf_2 fanout1217 (.A(net1218),
    .X(net1217));
 buf_2 fanout1218 (.A(_07281_),
    .X(net1218));
 buf_2 fanout1219 (.A(_07245_),
    .X(net1219));
 clkbuf_2 fanout1220 (.A(net1222),
    .X(net1220));
 clkbuf_2 fanout1221 (.A(net1222),
    .X(net1221));
 clkbuf_2 fanout1222 (.A(_05187_),
    .X(net1222));
 clkbuf_4 fanout1223 (.A(net1224),
    .X(net1223));
 buf_2 fanout1224 (.A(net1808),
    .X(net1224));
 clkbuf_4 fanout1225 (.A(_00169_),
    .X(net1225));
 buf_2 fanout1226 (.A(_00169_),
    .X(net1226));
 clkbuf_1 wire1227 (.A(net1228),
    .X(net1227));
 clkbuf_1 wire1228 (.A(_09171_),
    .X(net1228));
 buf_2 fanout1229 (.A(_07351_),
    .X(net1229));
 clkbuf_2 fanout1230 (.A(_07266_),
    .X(net1230));
 buf_2 fanout1231 (.A(_07262_),
    .X(net1231));
 buf_2 fanout1232 (.A(_07239_),
    .X(net1232));
 clkbuf_4 fanout1233 (.A(net1234),
    .X(net1233));
 clkbuf_4 fanout1234 (.A(net1235),
    .X(net1234));
 buf_2 fanout1235 (.A(net1651),
    .X(net1235));
 buf_2 fanout1236 (.A(net1238),
    .X(net1236));
 buf_2 fanout1237 (.A(net1238),
    .X(net1237));
 buf_2 fanout1238 (.A(_07068_),
    .X(net1238));
 clkbuf_4 fanout1239 (.A(net1240),
    .X(net1239));
 clkbuf_2 fanout1240 (.A(_07057_),
    .X(net1240));
 buf_2 fanout1241 (.A(net1717),
    .X(net1241));
 clkbuf_4 fanout1242 (.A(net1243),
    .X(net1242));
 buf_2 fanout1243 (.A(net1824),
    .X(net1243));
 clkbuf_4 fanout1244 (.A(net1649),
    .X(net1244));
 clkbuf_2 fanout1245 (.A(\digitop_pav2.access_inst.access_ctrl0.f_access_i ),
    .X(net1245));
 buf_2 fanout1246 (.A(net1248),
    .X(net1246));
 buf_1 fanout1247 (.A(net1248),
    .X(net1247));
 clkbuf_4 fanout1248 (.A(net1649),
    .X(net1248));
 buf_2 fanout1249 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.piex_dt_rx_done ),
    .X(net1249));
 buf_4 fanout1250 (.A(net1817),
    .X(net1250));
 clkbuf_4 fanout1251 (.A(\digitop_pav2.proc_ctrl_inst.cmdctr.cmdctr_end3 ),
    .X(net1251));
 buf_2 fanout1252 (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[4] ),
    .X(net1252));
 buf_2 fanout1253 (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[1] ),
    .X(net1253));
 buf_2 fanout1254 (.A(\digitop_pav2.proc_ctrl_inst.cmd.state[0] ),
    .X(net1254));
 clkbuf_4 fanout1255 (.A(net1259),
    .X(net1255));
 buf_2 fanout1256 (.A(net1258),
    .X(net1256));
 clkbuf_2 fanout1257 (.A(net1258),
    .X(net1257));
 clkbuf_4 fanout1258 (.A(net1707),
    .X(net1258));
 buf_2 fanout1259 (.A(net1706),
    .X(net1259));
 clkbuf_4 fanout1260 (.A(net1262),
    .X(net1260));
 buf_2 fanout1261 (.A(net1262),
    .X(net1261));
 buf_2 fanout1262 (.A(net1702),
    .X(net1262));
 buf_2 fanout1263 (.A(net1701),
    .X(net1263));
 clkbuf_4 fanout1264 (.A(net1266),
    .X(net1264));
 clkbuf_2 fanout1265 (.A(net1266),
    .X(net1265));
 buf_2 fanout1266 (.A(net1267),
    .X(net1266));
 clkbuf_2 fanout1267 (.A(net1658),
    .X(net1267));
 clkbuf_4 fanout1268 (.A(net1272),
    .X(net1268));
 clkbuf_4 fanout1269 (.A(net1272),
    .X(net1269));
 clkbuf_4 fanout1270 (.A(net1271),
    .X(net1270));
 clkbuf_2 fanout1271 (.A(net1272),
    .X(net1271));
 buf_2 fanout1272 (.A(net1691),
    .X(net1272));
 clkbuf_4 fanout1273 (.A(net1690),
    .X(net1273));
 clkbuf_2 fanout1274 (.A(net1689),
    .X(net1274));
 clkbuf_2 fanout1275 (.A(net1677),
    .X(net1275));
 buf_2 fanout1276 (.A(net1698),
    .X(net1276));
 clkbuf_2 fanout1277 (.A(net1681),
    .X(net1277));
 clkbuf_2 fanout1278 (.A(net1671),
    .X(net1278));
 clkbuf_2 fanout1279 (.A(net1669),
    .X(net1279));
 clkbuf_2 fanout1280 (.A(net1668),
    .X(net1280));
 clkbuf_2 fanout1281 (.A(net1674),
    .X(net1281));
 dlymetal6s2s_1 fanout1282 (.A(net1686),
    .X(net1282));
 clkbuf_4 fanout1283 (.A(net1285),
    .X(net1283));
 clkbuf_4 fanout1284 (.A(net1285),
    .X(net1284));
 buf_2 fanout1285 (.A(\digitop_pav2.fm0miller_inst.fm0x_ctrl.en_i ),
    .X(net1285));
 buf_2 fanout1286 (.A(net1288),
    .X(net1286));
 dlymetal6s2s_1 fanout1287 (.A(net1288),
    .X(net1287));
 clkbuf_2 fanout1288 (.A(net1289),
    .X(net1288));
 clkbuf_2 fanout1289 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[13] ),
    .X(net1289));
 clkbuf_4 fanout1290 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[7] ),
    .X(net1290));
 clkbuf_2 fanout1291 (.A(net1665),
    .X(net1291));
 clkbuf_2 fanout1292 (.A(net1293),
    .X(net1292));
 buf_2 fanout1293 (.A(net1662),
    .X(net1293));
 buf_2 fanout1294 (.A(net1295),
    .X(net1294));
 clkbuf_4 fanout1295 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[0] ),
    .X(net1295));
 clkbuf_4 fanout1296 (.A(_07041_),
    .X(net1296));
 buf_2 fanout1297 (.A(net1299),
    .X(net1297));
 buf_1 fanout1298 (.A(net1299),
    .X(net1298));
 buf_2 fanout1299 (.A(net1637),
    .X(net1299));
 buf_2 fanout1300 (.A(\digitop_pav2.pie_inst.fsm.pivot[6] ),
    .X(net1300));
 buf_2 fanout1301 (.A(\digitop_pav2.pie_inst.fsm.pivot[3] ),
    .X(net1301));
 buf_2 fanout1302 (.A(net1305),
    .X(net1302));
 buf_2 fanout1303 (.A(net1656),
    .X(net1303));
 clkbuf_4 fanout1304 (.A(net1305),
    .X(net1304));
 clkbuf_2 fanout1305 (.A(net1655),
    .X(net1305));
 buf_1 wire1306 (.A(_05419_),
    .X(net1306));
 clkbuf_4 fanout1307 (.A(_05525_),
    .X(net1307));
 clkbuf_2 fanout1308 (.A(_05525_),
    .X(net1308));
 buf_1 max_cap1309 (.A(_09501_),
    .X(net1309));
 clkbuf_2 fanout1310 (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.state[3] ),
    .X(net1310));
 buf_2 fanout1311 (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_fsm.en_pctr ),
    .X(net1311));
 clkbuf_4 fanout1312 (.A(_03660_),
    .X(net1312));
 clkbuf_2 fanout1313 (.A(_03660_),
    .X(net1313));
 buf_2 fanout1314 (.A(_11111_),
    .X(net1314));
 clkbuf_2 fanout1315 (.A(_11111_),
    .X(net1315));
 clkbuf_4 fanout1316 (.A(_07834_),
    .X(net1316));
 buf_2 fanout1317 (.A(_07834_),
    .X(net1317));
 clkbuf_4 fanout1318 (.A(_07418_),
    .X(net1318));
 clkbuf_4 fanout1319 (.A(_07417_),
    .X(net1319));
 buf_2 fanout1320 (.A(_10720_),
    .X(net1320));
 clkbuf_4 fanout1321 (.A(_10719_),
    .X(net1321));
 buf_6 fanout1322 (.A(net1829),
    .X(net1322));
 clkbuf_4 fanout1323 (.A(\digitop_pav2.access_inst.access_check0.fg_i[4] ),
    .X(net1323));
 buf_4 fanout1324 (.A(\digitop_pav2.access_inst.access_check0.fg_i[0] ),
    .X(net1324));
 buf_2 fanout1325 (.A(net1751),
    .X(net1325));
 buf_2 fanout1326 (.A(net1760),
    .X(net1326));
 clkbuf_4 fanout1327 (.A(net1329),
    .X(net1327));
 dlymetal6s2s_1 fanout1328 (.A(net1329),
    .X(net1328));
 clkbuf_2 fanout1329 (.A(net1344),
    .X(net1329));
 clkbuf_2 fanout1330 (.A(net1332),
    .X(net1330));
 clkbuf_2 fanout1331 (.A(net1332),
    .X(net1331));
 dlymetal6s2s_1 fanout1332 (.A(net1344),
    .X(net1332));
 clkbuf_2 fanout1333 (.A(net1334),
    .X(net1333));
 buf_1 fanout1334 (.A(net1344),
    .X(net1334));
 clkbuf_2 fanout1335 (.A(net1337),
    .X(net1335));
 clkbuf_2 fanout1336 (.A(net1337),
    .X(net1336));
 clkbuf_2 fanout1337 (.A(net1343),
    .X(net1337));
 clkbuf_2 fanout1338 (.A(net1339),
    .X(net1338));
 clkbuf_2 fanout1339 (.A(net1343),
    .X(net1339));
 clkbuf_2 fanout1340 (.A(net1342),
    .X(net1340));
 clkbuf_2 fanout1341 (.A(net1342),
    .X(net1341));
 buf_2 fanout1342 (.A(net1343),
    .X(net1342));
 clkbuf_2 fanout1343 (.A(net1344),
    .X(net1343));
 buf_2 fanout1344 (.A(\stadly_mpw03_erase_rise_9.Y ),
    .X(net1344));
 clkbuf_2 fanout1345 (.A(net1346),
    .X(net1345));
 clkbuf_2 fanout1346 (.A(net1350),
    .X(net1346));
 clkbuf_2 fanout1347 (.A(net1350),
    .X(net1347));
 buf_1 fanout1348 (.A(net1350),
    .X(net1348));
 clkbuf_2 fanout1349 (.A(net1350),
    .X(net1349));
 clkbuf_2 fanout1350 (.A(net1370),
    .X(net1350));
 clkbuf_2 fanout1351 (.A(net1355),
    .X(net1351));
 clkbuf_2 fanout1352 (.A(net1354),
    .X(net1352));
 clkbuf_2 fanout1353 (.A(net1354),
    .X(net1353));
 dlymetal6s2s_1 fanout1354 (.A(net1355),
    .X(net1354));
 dlymetal6s2s_1 fanout1355 (.A(net1370),
    .X(net1355));
 clkbuf_2 fanout1356 (.A(net1363),
    .X(net1356));
 buf_1 fanout1357 (.A(net1363),
    .X(net1357));
 clkbuf_2 fanout1358 (.A(net1363),
    .X(net1358));
 buf_1 fanout1359 (.A(net1363),
    .X(net1359));
 clkbuf_2 fanout1360 (.A(net1362),
    .X(net1360));
 clkbuf_2 fanout1361 (.A(net1362),
    .X(net1361));
 clkbuf_2 fanout1362 (.A(net1363),
    .X(net1362));
 clkbuf_2 fanout1363 (.A(net1370),
    .X(net1363));
 clkbuf_2 fanout1364 (.A(net1366),
    .X(net1364));
 clkbuf_2 fanout1365 (.A(net1366),
    .X(net1365));
 dlymetal6s2s_1 fanout1366 (.A(net1370),
    .X(net1366));
 clkbuf_2 fanout1367 (.A(net1369),
    .X(net1367));
 clkbuf_2 fanout1368 (.A(net1369),
    .X(net1368));
 clkbuf_2 fanout1369 (.A(net1370),
    .X(net1369));
 clkbuf_2 fanout1370 (.A(\stadly_mpw03_erase_rise_9.Y ),
    .X(net1370));
 clkbuf_2 fanout1371 (.A(net1372),
    .X(net1371));
 clkbuf_2 fanout1372 (.A(net1393),
    .X(net1372));
 clkbuf_2 fanout1373 (.A(net1375),
    .X(net1373));
 clkbuf_2 fanout1374 (.A(net1375),
    .X(net1374));
 clkbuf_2 fanout1375 (.A(net1393),
    .X(net1375));
 clkbuf_2 fanout1376 (.A(net1378),
    .X(net1376));
 clkbuf_2 fanout1377 (.A(net1378),
    .X(net1377));
 clkbuf_2 fanout1378 (.A(net1379),
    .X(net1378));
 clkbuf_2 fanout1379 (.A(net1393),
    .X(net1379));
 clkbuf_2 fanout1380 (.A(net1382),
    .X(net1380));
 clkbuf_2 fanout1381 (.A(net1382),
    .X(net1381));
 clkbuf_2 fanout1382 (.A(net1393),
    .X(net1382));
 clkbuf_2 fanout1383 (.A(net1385),
    .X(net1383));
 clkbuf_2 fanout1384 (.A(net1385),
    .X(net1384));
 clkbuf_2 fanout1385 (.A(net1393),
    .X(net1385));
 clkbuf_2 fanout1386 (.A(net1389),
    .X(net1386));
 clkbuf_2 fanout1387 (.A(net1389),
    .X(net1387));
 buf_1 fanout1388 (.A(net1389),
    .X(net1388));
 clkbuf_2 fanout1389 (.A(net1393),
    .X(net1389));
 clkbuf_2 fanout1390 (.A(net1392),
    .X(net1390));
 clkbuf_2 fanout1391 (.A(net1392),
    .X(net1391));
 clkbuf_2 fanout1392 (.A(net1393),
    .X(net1392));
 clkbuf_4 fanout1393 (.A(\stadly_mpw03_erase_rise_9.Y ),
    .X(net1393));
 buf_2 fanout1394 (.A(_03756_),
    .X(net1394));
 clkbuf_2 fanout1395 (.A(_03756_),
    .X(net1395));
 buf_2 fanout1396 (.A(net1397),
    .X(net1396));
 buf_2 fanout1397 (.A(_07060_),
    .X(net1397));
 clkbuf_4 fanout1398 (.A(net1399),
    .X(net1398));
 buf_2 fanout1399 (.A(_07060_),
    .X(net1399));
 clkbuf_4 fanout1400 (.A(_07060_),
    .X(net1400));
 clkbuf_4 fanout1401 (.A(net1402),
    .X(net1401));
 clkbuf_4 fanout1402 (.A(net1412),
    .X(net1402));
 clkbuf_4 fanout1403 (.A(net1404),
    .X(net1403));
 clkbuf_2 fanout1404 (.A(net1412),
    .X(net1404));
 clkbuf_4 fanout1405 (.A(net1408),
    .X(net1405));
 clkbuf_4 fanout1406 (.A(net1407),
    .X(net1406));
 clkbuf_4 fanout1407 (.A(net1408),
    .X(net1407));
 dlymetal6s2s_1 fanout1408 (.A(net1412),
    .X(net1408));
 clkbuf_4 fanout1409 (.A(net1410),
    .X(net1409));
 clkbuf_4 fanout1410 (.A(net1411),
    .X(net1410));
 buf_2 fanout1411 (.A(net1412),
    .X(net1411));
 clkbuf_4 fanout1412 (.A(net1413),
    .X(net1412));
 dlymetal6s2s_1 fanout1413 (.A(net1457),
    .X(net1413));
 clkbuf_4 fanout1414 (.A(net1418),
    .X(net1414));
 clkbuf_4 fanout1415 (.A(net1417),
    .X(net1415));
 clkbuf_4 fanout1416 (.A(net1417),
    .X(net1416));
 clkbuf_2 fanout1417 (.A(net1418),
    .X(net1417));
 clkbuf_2 fanout1418 (.A(net1421),
    .X(net1418));
 clkbuf_4 fanout1419 (.A(net1421),
    .X(net1419));
 buf_2 fanout1420 (.A(net1421),
    .X(net1420));
 buf_2 fanout1421 (.A(net1457),
    .X(net1421));
 clkbuf_4 fanout1422 (.A(net1423),
    .X(net1422));
 clkbuf_4 fanout1423 (.A(net1457),
    .X(net1423));
 clkbuf_4 fanout1424 (.A(net1427),
    .X(net1424));
 clkbuf_4 fanout1425 (.A(net1426),
    .X(net1425));
 buf_2 fanout1426 (.A(net1427),
    .X(net1426));
 clkbuf_2 fanout1427 (.A(net1436),
    .X(net1427));
 clkbuf_4 fanout1428 (.A(net1430),
    .X(net1428));
 buf_2 fanout1429 (.A(net1430),
    .X(net1429));
 clkbuf_2 fanout1430 (.A(net1436),
    .X(net1430));
 buf_2 fanout1431 (.A(net1433),
    .X(net1431));
 clkbuf_2 fanout1432 (.A(net1433),
    .X(net1432));
 clkbuf_4 fanout1433 (.A(net1436),
    .X(net1433));
 clkbuf_4 fanout1434 (.A(net1435),
    .X(net1434));
 buf_2 fanout1435 (.A(net1436),
    .X(net1435));
 clkbuf_4 fanout1436 (.A(net1457),
    .X(net1436));
 clkbuf_4 fanout1437 (.A(net1444),
    .X(net1437));
 clkbuf_2 fanout1438 (.A(net1443),
    .X(net1438));
 buf_2 fanout1439 (.A(net1440),
    .X(net1439));
 clkbuf_2 fanout1440 (.A(net1443),
    .X(net1440));
 clkbuf_4 fanout1441 (.A(net1443),
    .X(net1441));
 clkbuf_4 fanout1442 (.A(net1444),
    .X(net1442));
 clkbuf_2 fanout1443 (.A(net1444),
    .X(net1443));
 buf_2 fanout1444 (.A(net1704),
    .X(net1444));
 clkbuf_4 fanout1445 (.A(net1446),
    .X(net1445));
 clkbuf_4 fanout1446 (.A(net1456),
    .X(net1446));
 clkbuf_4 fanout1447 (.A(net1449),
    .X(net1447));
 clkbuf_4 fanout1448 (.A(net1449),
    .X(net1448));
 buf_2 fanout1449 (.A(net1456),
    .X(net1449));
 clkbuf_4 fanout1450 (.A(net1452),
    .X(net1450));
 buf_2 fanout1451 (.A(net1452),
    .X(net1451));
 clkbuf_2 fanout1452 (.A(net1453),
    .X(net1452));
 clkbuf_2 fanout1453 (.A(net1456),
    .X(net1453));
 clkbuf_4 fanout1454 (.A(net1456),
    .X(net1454));
 clkbuf_2 fanout1455 (.A(net1456),
    .X(net1455));
 clkbuf_4 fanout1456 (.A(net1704),
    .X(net1456));
 clkbuf_8 fanout1457 (.A(net1703),
    .X(net1457));
 buf_2 fanout1458 (.A(_03839_),
    .X(net1458));
 dlymetal6s2s_1 fanout1459 (.A(_03839_),
    .X(net1459));
 buf_2 fanout1460 (.A(_03754_),
    .X(net1460));
 clkbuf_2 fanout1461 (.A(_03754_),
    .X(net1461));
 buf_2 fanout1462 (.A(net1463),
    .X(net1462));
 clkbuf_2 fanout1463 (.A(_03753_),
    .X(net1463));
 clkbuf_2 max_cap1464 (.A(_09630_),
    .X(net1464));
 clkbuf_1 max_cap1465 (.A(_09619_),
    .X(net1465));
 buf_1 max_cap1466 (.A(_09591_),
    .X(net1466));
 buf_2 fanout1467 (.A(_03826_),
    .X(net1467));
 buf_2 fanout1468 (.A(_03782_),
    .X(net1468));
 clkbuf_2 fanout1469 (.A(_03782_),
    .X(net1469));
 buf_2 fanout1470 (.A(_03758_),
    .X(net1470));
 buf_2 fanout1471 (.A(net1472),
    .X(net1471));
 clkbuf_4 fanout1472 (.A(_03757_),
    .X(net1472));
 buf_1 max_cap1473 (.A(_03731_),
    .X(net1473));
 clkbuf_2 fanout1474 (.A(net1475),
    .X(net1474));
 dlymetal6s2s_1 fanout1475 (.A(net1476),
    .X(net1475));
 clkbuf_2 fanout1476 (.A(_07113_),
    .X(net1476));
 clkbuf_4 fanout1477 (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[4] ),
    .X(net1477));
 buf_2 fanout1478 (.A(net1479),
    .X(net1478));
 clkbuf_2 fanout1479 (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_iface.addr_ff[3] ),
    .X(net1479));
 buf_2 fanout1480 (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rd_end_i ),
    .X(net1480));
 buf_4 fanout1481 (.A(\digitop_pav2.testctrl_pav2.inst_mbform.inst_type.tm_mbist_i ),
    .X(net1481));
 buf_2 fanout1482 (.A(net1483),
    .X(net1482));
 clkbuf_4 fanout1483 (.A(\digitop_pav2.cal_inst.calx_mux.en_calx_test_i ),
    .X(net1483));
 buf_2 fanout1484 (.A(\digitop_pav2.testctrl_pav2.inst_mode.state[4] ),
    .X(net1484));
 buf_1 fanout1485 (.A(\digitop_pav2.testctrl_pav2.inst_mode.state[4] ),
    .X(net1485));
 buf_2 fanout1486 (.A(\digitop_pav2.testctrl_pav2.inst_mode.state[3] ),
    .X(net1486));
 clkbuf_2 fanout1487 (.A(\digitop_pav2.testctrl_pav2.inst_mode.state[2] ),
    .X(net1487));
 buf_1 fanout1488 (.A(\digitop_pav2.testctrl_pav2.inst_mode.state[2] ),
    .X(net1488));
 clkbuf_2 fanout1489 (.A(\digitop_pav2.testctrl_pav2.inst_mode.state[1] ),
    .X(net1489));
 buf_2 fanout1490 (.A(\digitop_pav2.testctrl_pav2.inst_mode.state[0] ),
    .X(net1490));
 buf_1 fanout1491 (.A(\digitop_pav2.testctrl_pav2.inst_mode.state[0] ),
    .X(net1491));
 clkbuf_4 fanout1492 (.A(net1500),
    .X(net1492));
 buf_2 fanout1493 (.A(net1494),
    .X(net1493));
 buf_4 fanout1494 (.A(net1500),
    .X(net1494));
 buf_4 fanout1495 (.A(net1498),
    .X(net1495));
 buf_2 fanout1496 (.A(net1498),
    .X(net1496));
 buf_4 fanout1497 (.A(net1498),
    .X(net1497));
 buf_2 fanout1498 (.A(net1500),
    .X(net1498));
 buf_4 fanout1499 (.A(net1500),
    .X(net1499));
 buf_2 fanout1500 (.A(_07166_),
    .X(net1500));
 buf_2 fanout1501 (.A(net1502),
    .X(net1501));
 clkbuf_2 fanout1502 (.A(net1503),
    .X(net1502));
 clkbuf_4 fanout1503 (.A(net69),
    .X(net1503));
 buf_2 fanout1504 (.A(net67),
    .X(net1504));
 clkbuf_4 fanout1505 (.A(net1575),
    .X(net1505));
 clkbuf_4 fanout1506 (.A(net1514),
    .X(net1506));
 buf_2 fanout1507 (.A(net1514),
    .X(net1507));
 clkbuf_4 fanout1508 (.A(net1514),
    .X(net1508));
 clkbuf_2 fanout1509 (.A(net1514),
    .X(net1509));
 clkbuf_4 fanout1510 (.A(net1511),
    .X(net1510));
 buf_2 fanout1511 (.A(net1513),
    .X(net1511));
 clkbuf_4 fanout1512 (.A(net1513),
    .X(net1512));
 clkbuf_2 fanout1513 (.A(net1514),
    .X(net1513));
 clkbuf_2 fanout1514 (.A(net1575),
    .X(net1514));
 clkbuf_4 fanout1515 (.A(net1517),
    .X(net1515));
 clkbuf_2 fanout1516 (.A(net1517),
    .X(net1516));
 clkbuf_4 fanout1517 (.A(net1518),
    .X(net1517));
 buf_2 fanout1518 (.A(net1575),
    .X(net1518));
 clkbuf_4 fanout1519 (.A(net1521),
    .X(net1519));
 clkbuf_4 fanout1520 (.A(net1521),
    .X(net1520));
 clkbuf_4 fanout1521 (.A(net1548),
    .X(net1521));
 clkbuf_4 fanout1522 (.A(net1525),
    .X(net1522));
 clkbuf_2 fanout1523 (.A(net1525),
    .X(net1523));
 clkbuf_4 fanout1524 (.A(net1525),
    .X(net1524));
 buf_2 fanout1525 (.A(net1548),
    .X(net1525));
 clkbuf_4 fanout1526 (.A(net1530),
    .X(net1526));
 clkbuf_2 fanout1527 (.A(net1530),
    .X(net1527));
 clkbuf_4 fanout1528 (.A(net1530),
    .X(net1528));
 clkbuf_4 fanout1529 (.A(net1530),
    .X(net1529));
 buf_2 fanout1530 (.A(net1548),
    .X(net1530));
 clkbuf_4 fanout1531 (.A(net1534),
    .X(net1531));
 buf_2 fanout1532 (.A(net1534),
    .X(net1532));
 clkbuf_4 fanout1533 (.A(net1534),
    .X(net1533));
 buf_2 fanout1534 (.A(net1539),
    .X(net1534));
 clkbuf_4 fanout1535 (.A(net1539),
    .X(net1535));
 buf_2 fanout1536 (.A(net1539),
    .X(net1536));
 clkbuf_4 fanout1537 (.A(net1539),
    .X(net1537));
 clkbuf_2 fanout1538 (.A(net1539),
    .X(net1538));
 clkbuf_2 fanout1539 (.A(net1548),
    .X(net1539));
 clkbuf_4 fanout1540 (.A(net1542),
    .X(net1540));
 clkbuf_4 fanout1541 (.A(net1542),
    .X(net1541));
 buf_2 fanout1542 (.A(net1547),
    .X(net1542));
 clkbuf_4 fanout1543 (.A(net1547),
    .X(net1543));
 clkbuf_2 fanout1544 (.A(net1547),
    .X(net1544));
 clkbuf_4 fanout1545 (.A(net1547),
    .X(net1545));
 clkbuf_2 fanout1546 (.A(net1547),
    .X(net1546));
 clkbuf_2 fanout1547 (.A(net1548),
    .X(net1547));
 buf_2 fanout1548 (.A(net1575),
    .X(net1548));
 clkbuf_4 fanout1549 (.A(net1552),
    .X(net1549));
 clkbuf_2 fanout1550 (.A(net1552),
    .X(net1550));
 clkbuf_4 fanout1551 (.A(net1552),
    .X(net1551));
 clkbuf_2 fanout1552 (.A(net1553),
    .X(net1552));
 clkbuf_4 fanout1553 (.A(net1574),
    .X(net1553));
 clkbuf_4 fanout1554 (.A(net1574),
    .X(net1554));
 buf_2 fanout1555 (.A(net1574),
    .X(net1555));
 clkbuf_4 fanout1556 (.A(net1559),
    .X(net1556));
 clkbuf_2 fanout1557 (.A(net1559),
    .X(net1557));
 clkbuf_4 fanout1558 (.A(net1559),
    .X(net1558));
 buf_2 fanout1559 (.A(net1564),
    .X(net1559));
 clkbuf_4 fanout1560 (.A(net1564),
    .X(net1560));
 clkbuf_2 fanout1561 (.A(net1564),
    .X(net1561));
 clkbuf_4 fanout1562 (.A(net1564),
    .X(net1562));
 buf_2 fanout1563 (.A(net1564),
    .X(net1563));
 clkbuf_2 fanout1564 (.A(net1574),
    .X(net1564));
 clkbuf_4 fanout1565 (.A(net1568),
    .X(net1565));
 clkbuf_2 fanout1566 (.A(net1568),
    .X(net1566));
 clkbuf_4 fanout1567 (.A(net1568),
    .X(net1567));
 buf_2 fanout1568 (.A(net1573),
    .X(net1568));
 clkbuf_4 fanout1569 (.A(net1573),
    .X(net1569));
 clkbuf_2 fanout1570 (.A(net1573),
    .X(net1570));
 clkbuf_4 fanout1571 (.A(net1573),
    .X(net1571));
 clkbuf_2 fanout1572 (.A(net1573),
    .X(net1572));
 clkbuf_2 fanout1573 (.A(net1574),
    .X(net1573));
 buf_2 fanout1574 (.A(net1575),
    .X(net1574));
 clkbuf_4 fanout1575 (.A(net66),
    .X(net1575));
 clkbuf_4 fanout1576 (.A(net1578),
    .X(net1576));
 clkbuf_2 fanout1577 (.A(net1578),
    .X(net1577));
 buf_2 fanout1578 (.A(net1581),
    .X(net1578));
 clkbuf_4 fanout1579 (.A(net1580),
    .X(net1579));
 clkbuf_4 fanout1580 (.A(net1581),
    .X(net1580));
 buf_2 fanout1581 (.A(net66),
    .X(net1581));
 conb_1 _24114__1582 (.LO(net1582));
 conb_1 \digitop_pav2.fm0miller_inst.fm0x_tx.muxdata_fmdata_1_1609  (.LO(net1609));
 conb_1 \digitop_pav2.fm0miller_inst.fm0x_tx.muxdata_fmdata_1_1616  (.HI(net1616));
 dlygate4sd3_1 hold2 (.A(net1623),
    .X(net1618));
 dlygate4sd3_1 hold3 (.A(\digitop_pav2.g_auth_obu ),
    .X(net1619));
 dlygate4sd3_1 hold4 (.A(net1008),
    .X(net1620));
 dlygate4sd3_1 hold5 (.A(net1007),
    .X(net1621));
 dlygate4sd3_1 hold6 (.A(net1633),
    .X(net1622));
 dlygate4sd3_1 hold7 (.A(net1627),
    .X(net1623));
 dlygate4sd3_1 hold8 (.A(net1618),
    .X(net1624));
 dlygate4sd3_1 hold9 (.A(net1630),
    .X(net1625));
 dlygate4sd3_1 hold10 (.A(net1617),
    .X(net1626));
 dlygate4sd3_1 hold11 (.A(_07851_),
    .X(net1627));
 dlygate4sd3_1 hold12 (.A(net1632),
    .X(net1628));
 dlygate4sd3_1 hold13 (.A(net1622),
    .X(net1629));
 dlygate4sd3_1 hold14 (.A(\digitop_pav2.proc_ctrl_inst.cmd.g_sec_auth_o ),
    .X(net1630));
 dlygate4sd3_1 hold15 (.A(net1625),
    .X(net1631));
 dlygate4sd3_1 hold16 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.cmdfsm_cgen.en_g_sec_i ),
    .X(net1632));
 dlygate4sd3_1 hold17 (.A(net1628),
    .X(net1633));
 dlygate4sd3_1 hold18 (.A(\digitop_pav2.memctrl_inst.busy_ff ),
    .X(net1634));
 dlygate4sd3_1 hold19 (.A(\digitop_pav2.access_inst.access_ctrl0.nvm_busy_i ),
    .X(net1635));
 dlygate4sd3_1 hold20 (.A(_09653_),
    .X(net1636));
 dlygate4sd3_1 hold21 (.A(\digitop_pav2.crc_inst.dt_rx_i ),
    .X(net1637));
 dlygate4sd3_1 hold22 (.A(net1299),
    .X(net1638));
 dlygate4sd3_1 hold23 (.A(net1657),
    .X(net1639));
 dlygate4sd3_1 hold24 (.A(net817),
    .X(net1640));
 dlygate4sd3_1 hold25 (.A(net813),
    .X(net1641));
 dlygate4sd3_1 hold26 (.A(_00680_),
    .X(net1642));
 dlygate4sd3_1 hold27 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[8] ),
    .X(net1643));
 dlygate4sd3_1 hold28 (.A(_07327_),
    .X(net1644));
 dlygate4sd3_1 hold29 (.A(net1661),
    .X(net1645));
 dlygate4sd3_1 hold30 (.A(net819),
    .X(net1646));
 dlygate4sd3_1 hold31 (.A(_03706_),
    .X(net1647));
 dlygate4sd3_1 hold32 (.A(_00495_),
    .X(net1648));
 dlygate4sd3_1 hold33 (.A(net1667),
    .X(net1649));
 dlygate4sd3_1 hold34 (.A(net1244),
    .X(net1650));
 dlygate4sd3_1 hold35 (.A(_07086_),
    .X(net1651));
 dlygate4sd3_1 hold36 (.A(net1235),
    .X(net1652));
 dlygate4sd3_1 hold37 (.A(_03705_),
    .X(net1653));
 dlygate4sd3_1 hold38 (.A(_00896_),
    .X(net1654));
 dlygate4sd3_1 hold39 (.A(\digitop_pav2.crc_inst.dt_rx_en_i ),
    .X(net1655));
 dlygate4sd3_1 hold40 (.A(net1305),
    .X(net1656));
 dlygate4sd3_1 hold41 (.A(_07380_),
    .X(net1657));
 dlygate4sd3_1 hold42 (.A(\digitop_pav2.ack_inst.g_ack_i ),
    .X(net1658));
 dlygate4sd3_1 hold43 (.A(_07325_),
    .X(net1659));
 dlygate4sd3_1 hold44 (.A(_07326_),
    .X(net1660));
 dlygate4sd3_1 hold45 (.A(_07335_),
    .X(net1661));
 dlygate4sd3_1 hold46 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[2] ),
    .X(net1662));
 dlygate4sd3_1 hold47 (.A(_07279_),
    .X(net1663));
 dlygate4sd3_1 hold48 (.A(_07333_),
    .X(net1664));
 dlygate4sd3_1 hold49 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[6] ),
    .X(net1665));
 dlygate4sd3_1 hold50 (.A(_07283_),
    .X(net1666));
 dlygate4sd3_1 hold51 (.A(\digitop_pav2.access_inst.access_ctrl0.f_access_i ),
    .X(net1667));
 dlygate4sd3_1 hold52 (.A(net1683),
    .X(net1668));
 dlygate4sd3_1 hold53 (.A(net1280),
    .X(net1669));
 dlygate4sd3_1 hold54 (.A(_00275_),
    .X(net1670));
 dlygate4sd3_1 hold55 (.A(net1680),
    .X(net1671));
 dlygate4sd3_1 hold56 (.A(net1278),
    .X(net1672));
 dlygate4sd3_1 hold57 (.A(_00270_),
    .X(net1673));
 dlygate4sd3_1 hold58 (.A(net1685),
    .X(net1674));
 dlygate4sd3_1 hold59 (.A(net1281),
    .X(net1675));
 dlygate4sd3_1 hold60 (.A(_00350_),
    .X(net1676));
 dlygate4sd3_1 hold61 (.A(net1688),
    .X(net1677));
 dlygate4sd3_1 hold62 (.A(net1275),
    .X(net1678));
 dlygate4sd3_1 hold63 (.A(_00268_),
    .X(net1679));
 dlygate4sd3_1 hold64 (.A(\digitop_pav2.g_queryadj ),
    .X(net1680));
 dlygate4sd3_1 hold65 (.A(net1671),
    .X(net1681));
 dlygate4sd3_1 hold66 (.A(_00271_),
    .X(net1682));
 dlygate4sd3_1 hold67 (.A(\digitop_pav2.g_queryrep ),
    .X(net1683));
 dlygate4sd3_1 hold68 (.A(_00351_),
    .X(net1684));
 dlygate4sd3_1 hold69 (.A(\digitop_pav2.g_reqrn ),
    .X(net1685));
 dlygate4sd3_1 hold70 (.A(net1674),
    .X(net1686));
 dlygate4sd3_1 hold71 (.A(_00349_),
    .X(net1687));
 dlygate4sd3_1 hold72 (.A(\digitop_pav2.g_query ),
    .X(net1688));
 dlygate4sd3_1 hold73 (.A(net1677),
    .X(net1689));
 dlygate4sd3_1 hold74 (.A(net1693),
    .X(net1690));
 dlygate4sd3_1 hold75 (.A(net1273),
    .X(net1691));
 dlygate4sd3_1 hold76 (.A(_00168_),
    .X(net1692));
 dlygate4sd3_1 hold77 (.A(\digitop_pav2.g_select ),
    .X(net1693));
 dlygate4sd3_1 hold78 (.A(net1708),
    .X(net1694));
 dlygate4sd3_1 hold79 (.A(_07069_),
    .X(net1695));
 dlygate4sd3_1 hold80 (.A(_07322_),
    .X(net1696));
 dlygate4sd3_1 hold81 (.A(net1214),
    .X(net1697));
 dlygate4sd3_1 hold82 (.A(net1709),
    .X(net1698));
 dlygate4sd3_1 hold83 (.A(net1276),
    .X(net1699));
 dlygate4sd3_1 hold84 (.A(_07320_),
    .X(net1700));
 dlygate4sd3_1 hold85 (.A(\digitop_pav2.access_inst.access_check0.g_read_i ),
    .X(net1701));
 dlygate4sd3_1 hold86 (.A(net1263),
    .X(net1702));
 dlygate4sd3_1 hold87 (.A(\digitop_pav2.aes128_inst.aes128_counter.rst_b_i ),
    .X(net1703));
 dlygate4sd3_1 hold88 (.A(net1457),
    .X(net1704));
 dlygate4sd3_1 hold89 (.A(\digitop_pav2.glue_inst.mbus_rd_en_o ),
    .X(net1705));
 dlygate4sd3_1 hold90 (.A(\digitop_pav2.access_inst.access_check0.g_activate_i ),
    .X(net1706));
 dlygate4sd3_1 hold91 (.A(net1259),
    .X(net1707));
 dlygate4sd3_1 hold92 (.A(\digitop_pav2.access_inst.access_check0.g_propwrite_i ),
    .X(net1708));
 dlygate4sd3_1 hold93 (.A(\digitop_pav2.access_inst.access_check0.g_write_i ),
    .X(net1709));
 dlygate4sd3_1 hold94 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[11] ),
    .X(net1710));
 dlygate4sd3_1 hold95 (.A(_07359_),
    .X(net1711));
 dlygate4sd3_1 hold96 (.A(_07368_),
    .X(net1712));
 dlygate4sd3_1 hold97 (.A(net1724),
    .X(net1713));
 dlygate4sd3_1 hold98 (.A(_10696_),
    .X(net1714));
 dlygate4sd3_1 hold99 (.A(_10702_),
    .X(net1715));
 dlygate4sd3_1 hold100 (.A(_10712_),
    .X(net1716));
 dlygate4sd3_1 hold101 (.A(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[0] ),
    .X(net1717));
 dlygate4sd3_1 hold102 (.A(net1241),
    .X(net1718));
 dlygate4sd3_1 hold103 (.A(_10697_),
    .X(net1719));
 dlygate4sd3_1 hold104 (.A(_10700_),
    .X(net1720));
 dlygate4sd3_1 hold105 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.state[1] ),
    .X(net1721));
 dlygate4sd3_1 hold106 (.A(net1723),
    .X(net1722));
 dlygate4sd3_1 hold107 (.A(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[2] ),
    .X(net1723));
 dlygate4sd3_1 hold108 (.A(\digitop_pav2.proc_ctrl_inst.cmd.state_pro_i[1] ),
    .X(net1724));
 dlygate4sd3_1 hold109 (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.dis_blf_fc_b ),
    .X(net1725));
 dlygate4sd3_1 hold110 (.A(_00210_),
    .X(net1726));
 dlygate4sd3_1 hold111 (.A(\digitop_pav2.proc_ctrl_inst.timeout.ctr.pass_t2 ),
    .X(net1727));
 dlygate4sd3_1 hold112 (.A(\digitop_pav2.pass_t2 ),
    .X(net1728));
 dlygate4sd3_1 hold113 (.A(\digitop_pav2.access_inst.access_transceiver0.handle_i[15] ),
    .X(net1729));
 dlygate4sd3_1 hold114 (.A(_07443_),
    .X(net1730));
 dlygate4sd3_1 hold115 (.A(_07444_),
    .X(net1731));
 dlygate4sd3_1 hold116 (.A(\digitop_pav2.func_rng_data[7] ),
    .X(net1732));
 dlygate4sd3_1 hold117 (.A(_05138_),
    .X(net1733));
 dlygate4sd3_1 hold118 (.A(\digitop_pav2.func_rng_data[1] ),
    .X(net1734));
 dlygate4sd3_1 hold119 (.A(_08889_),
    .X(net1735));
 dlygate4sd3_1 hold120 (.A(\digitop_pav2.func_rng_data[0] ),
    .X(net1736));
 dlygate4sd3_1 hold121 (.A(_08877_),
    .X(net1737));
 dlygate4sd3_1 hold122 (.A(\digitop_pav2.memctrl_inst.extra_dt_i[13] ),
    .X(net1738));
 dlygate4sd3_1 hold123 (.A(_05003_),
    .X(net1739));
 dlygate4sd3_1 hold124 (.A(_05008_),
    .X(net1740));
 dlygate4sd3_1 hold125 (.A(\digitop_pav2.func_rng_data[3] ),
    .X(net1741));
 dlygate4sd3_1 hold126 (.A(_08887_),
    .X(net1742));
 dlygate4sd3_1 hold127 (.A(\digitop_pav2.memctrl_inst.extra_dt_i[14] ),
    .X(net1743));
 dlygate4sd3_1 hold128 (.A(_05009_),
    .X(net1744));
 dlygate4sd3_1 hold129 (.A(_05015_),
    .X(net1745));
 dlygate4sd3_1 hold130 (.A(\digitop_pav2.memctrl_inst.extra_dt_i[12] ),
    .X(net1746));
 dlygate4sd3_1 hold131 (.A(_04995_),
    .X(net1747));
 dlygate4sd3_1 hold132 (.A(_05001_),
    .X(net1748));
 dlygate4sd3_1 hold133 (.A(\digitop_pav2.memctrl_inst.extra_dt_i[15] ),
    .X(net1749));
 dlygate4sd3_1 hold134 (.A(_05022_),
    .X(net1750));
 dlygate4sd3_1 hold135 (.A(\digitop_pav2.boot_inst.boot_proc0.proc_stage[1] ),
    .X(net1751));
 dlygate4sd3_1 hold136 (.A(net1325),
    .X(net1752));
 dlygate4sd3_1 hold137 (.A(_07918_),
    .X(net1753));
 dlygate4sd3_1 hold138 (.A(_04814_),
    .X(net1754));
 dlygate4sd3_1 hold139 (.A(\digitop_pav2.boot_inst.boot_ctrl0.ctrl_crc_en ),
    .X(net1755));
 dlygate4sd3_1 hold140 (.A(_07885_),
    .X(net1756));
 dlygate4sd3_1 hold141 (.A(_07886_),
    .X(net1757));
 dlygate4sd3_1 hold142 (.A(_07896_),
    .X(net1758));
 dlygate4sd3_1 hold143 (.A(_04815_),
    .X(net1759));
 dlygate4sd3_1 hold144 (.A(\digitop_pav2.boot_inst.boot_proc0.proc_stage[0] ),
    .X(net1760));
 dlygate4sd3_1 hold145 (.A(net1326),
    .X(net1761));
 dlygate4sd3_1 hold146 (.A(_07911_),
    .X(net1762));
 dlygate4sd3_1 hold147 (.A(_07912_),
    .X(net1763));
 dlygate4sd3_1 hold148 (.A(_07928_),
    .X(net1764));
 dlygate4sd3_1 hold149 (.A(\digitop_pav2.func_rng_data[4] ),
    .X(net1765));
 dlygate4sd3_1 hold150 (.A(\digitop_pav2.func_rng_data[2] ),
    .X(net1766));
 dlygate4sd3_1 hold151 (.A(\digitop_pav2.func_rng_data[10] ),
    .X(net1767));
 dlygate4sd3_1 hold152 (.A(\digitop_pav2.func_rng_data[6] ),
    .X(net1768));
 dlygate4sd3_1 hold153 (.A(\digitop_pav2.func_rng_data[12] ),
    .X(net1769));
 dlygate4sd3_1 hold154 (.A(\digitop_pav2.func_rng_data[5] ),
    .X(net1770));
 dlygate4sd3_1 hold155 (.A(\digitop_pav2.boot_inst.boot_ctrl0.proc_boot_end_i ),
    .X(net1771));
 dlygate4sd3_1 hold156 (.A(_07838_),
    .X(net1772));
 dlygate4sd3_1 hold157 (.A(_07842_),
    .X(net1773));
 dlygate4sd3_1 hold158 (.A(_07919_),
    .X(net1774));
 dlygate4sd3_1 hold159 (.A(_04817_),
    .X(net1775));
 dlygate4sd3_1 hold160 (.A(\digitop_pav2.func_rng_data[14] ),
    .X(net1776));
 dlygate4sd3_1 hold161 (.A(\digitop_pav2.boot_inst.boot_ctrl0.prev_busy ),
    .X(net1777));
 dlygate4sd3_1 hold162 (.A(_07840_),
    .X(net1778));
 dlygate4sd3_1 hold163 (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[0] ),
    .X(net1779));
 dlygate4sd3_1 hold164 (.A(\digitop_pav2.func_rng_data[9] ),
    .X(net1780));
 dlygate4sd3_1 hold165 (.A(\digitop_pav2.func_rng_data[13] ),
    .X(net1781));
 dlygate4sd3_1 hold166 (.A(\digitop_pav2.func_rng_data[8] ),
    .X(net1782));
 dlygate4sd3_1 hold167 (.A(\digitop_pav2.boot_inst.boot_ctrl0.replay ),
    .X(net1783));
 dlygate4sd3_1 hold168 (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[7] ),
    .X(net1784));
 dlygate4sd3_1 hold169 (.A(_11119_),
    .X(net1785));
 dlygate4sd3_1 hold170 (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[15] ),
    .X(net1786));
 dlygate4sd3_1 hold171 (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[8] ),
    .X(net1787));
 dlygate4sd3_1 hold172 (.A(\digitop_pav2.access_inst.access_check0.fg_i[13] ),
    .X(net1788));
 dlygate4sd3_1 hold173 (.A(\digitop_pav2.stadly_memctrl_wr_dt14_0.A ),
    .X(net1789));
 dlygate4sd3_1 hold174 (.A(\digitop_pav2.access_inst.access_check0.fg_i[11] ),
    .X(net1790));
 dlygate4sd3_1 hold175 (.A(\digitop_pav2.stadly_memctrl_wr_dt12_0.A ),
    .X(net1791));
 dlygate4sd3_1 hold176 (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[10] ),
    .X(net1792));
 dlygate4sd3_1 hold177 (.A(\digitop_pav2.stadly_memctrl_wr_dt10_0.A ),
    .X(net1793));
 dlygate4sd3_1 hold178 (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[6] ),
    .X(net1794));
 dlygate4sd3_1 hold179 (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[9] ),
    .X(net1795));
 dlygate4sd3_1 hold180 (.A(\digitop_pav2.stadly_memctrl_wr_dt9_0.A ),
    .X(net1796));
 dlygate4sd3_1 hold181 (.A(\digitop_pav2.access_inst.access_check0.fg_i[10] ),
    .X(net1797));
 dlygate4sd3_1 hold182 (.A(\digitop_pav2.stadly_memctrl_wr_dt11_0.A ),
    .X(net1798));
 dlygate4sd3_1 hold183 (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[4] ),
    .X(net1799));
 dlygate4sd3_1 hold184 (.A(\digitop_pav2.stadly_memctrl_wr_dt4_0.A ),
    .X(net1800));
 dlygate4sd3_1 hold185 (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[3] ),
    .X(net1801));
 dlygate4sd3_1 hold186 (.A(\digitop_pav2.stadly_memctrl_wr_dt3_0.A ),
    .X(net1802));
 dlygate4sd3_1 hold187 (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[13] ),
    .X(net1803));
 dlygate4sd3_1 hold188 (.A(\digitop_pav2.boot_inst.boot_proc0.boot_crc16_prl0.crc16[2] ),
    .X(net1804));
 dlygate4sd3_1 hold189 (.A(\digitop_pav2.stadly_memctrl_wr_dt2_0.A ),
    .X(net1805));
 dlygate4sd3_1 hold190 (.A(\digitop_pav2.func_rng_data[11] ),
    .X(net1806));
 dlygate4sd3_1 hold191 (.A(\digitop_pav2.pie_inst.delend_o ),
    .X(net1807));
 dlygate4sd3_1 hold192 (.A(\digitop_pav2.proc_ctrl_inst.cmd.rst_b_i ),
    .X(net1808));
 dlygate4sd3_1 hold193 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.ebv_rst_b ),
    .X(net1809));
 dlygate4sd3_1 hold194 (.A(ff_prog_ff),
    .X(net1810));
 dlygate4sd3_1 hold195 (.A(s2_rst_ff),
    .X(net1811));
 dlygate4sd3_1 hold196 (.A(s3_rst_ff),
    .X(net1812));
 dlygate4sd3_1 hold197 (.A(s3_set_ff),
    .X(net1813));
 dlygate4sd3_1 hold198 (.A(sl_rst_ff),
    .X(net1814));
 dlygate4sd3_1 hold199 (.A(ff_erase_ff),
    .X(net1815));
 dlygate4sd3_1 hold200 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.mode ),
    .X(net1816));
 dlygate4sd3_1 hold201 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.mode ),
    .X(net1817));
 dlygate4sd3_1 hold202 (.A(s2_set_ff),
    .X(net1818));
 dlygate4sd3_1 hold203 (.A(s1_set_ff),
    .X(net1819));
 dlygate4sd3_1 hold204 (.A(s1_rst_ff),
    .X(net1820));
 dlygate4sd3_1 hold205 (.A(sl_set_ff),
    .X(net1821));
 dlygate4sd3_1 hold206 (.A(ff_prog_ff2),
    .X(net1822));
 dlygate4sd3_1 hold207 (.A(ff_erase_ff2),
    .X(net1823));
 dlygate4sd3_1 hold208 (.A(\digitop_pav2.proc_ctrl_inst.cmdfsm.rn_rst_b ),
    .X(net1824));
 dlygate4sd3_1 hold209 (.A(\digitop_pav2.sync_inst.inst_rstx.sync_rstx_DONT_TOUCH.genblk1.genblk1[0].sync_pav2_clkx_delay_DONT_TOUCH.A ),
    .X(net1825));
 dlygate4sd3_1 hold210 (.A(\digitop_pav2.cal_inst.dtest.calx_dtest_clk.ref_pulse_sync_o ),
    .X(net1826));
 dlygate4sd3_1 hold211 (.A(\digitop_pav2.sync_inst.inst_clkx.inst_rngx.inst_pup_en.pup_ctr[5] ),
    .X(net1827));
 dlygate4sd3_1 hold212 (.A(_11104_),
    .X(net1828));
 dlygate4sd3_1 hold213 (.A(\digitop_pav2.access_inst.access_check0.permalock_tid_i ),
    .X(net1829));
 dlygate4sd3_1 hold214 (.A(s3_rst_ff2),
    .X(net1830));
 dlygate4sd3_1 hold215 (.A(_00355_),
    .X(net1831));
 dlygate4sd3_1 hold216 (.A(\digitop_pav2.sync_inst.inst_clkx.inst_blf.inst_en.pass_t2_ff ),
    .X(net1832));
 dlygate4sd3_1 hold217 (.A(s2_rst_ff2),
    .X(net1833));
 dlygate4sd3_1 hold218 (.A(_00356_),
    .X(net1834));
 dlygate4sd3_1 hold219 (.A(sl_rst_ff2),
    .X(net1835));
 dlygate4sd3_1 hold220 (.A(_00354_),
    .X(net1836));
 dlygate4sd3_1 hold221 (.A(s1_rst_ff2),
    .X(net1837));
 dlygate4sd3_1 hold222 (.A(_00489_),
    .X(net1838));
 dlygate4sd3_1 hold223 (.A(\digitop_pav2.sync_inst.inst_rstx.trigger_DONT_TOUCH1.Q ),
    .X(net1839));
 diode_2 ANTENNA_1 (.DIODE(_02192_));
 diode_2 ANTENNA_2 (.DIODE(_02192_));
 diode_2 ANTENNA_3 (.DIODE(_02192_));
 diode_2 ANTENNA_4 (.DIODE(_02192_));
 diode_2 ANTENNA_5 (.DIODE(_02826_));
 diode_2 ANTENNA_6 (.DIODE(_03254_));
 diode_2 ANTENNA_7 (.DIODE(_03766_));
 diode_2 ANTENNA_8 (.DIODE(_03808_));
 diode_2 ANTENNA_9 (.DIODE(_03824_));
 diode_2 ANTENNA_10 (.DIODE(_03891_));
 diode_2 ANTENNA_11 (.DIODE(_04189_));
 diode_2 ANTENNA_12 (.DIODE(_04189_));
 diode_2 ANTENNA_13 (.DIODE(_05019_));
 diode_2 ANTENNA_14 (.DIODE(_05572_));
 diode_2 ANTENNA_15 (.DIODE(_05621_));
 diode_2 ANTENNA_16 (.DIODE(_06411_));
 diode_2 ANTENNA_17 (.DIODE(_06411_));
 diode_2 ANTENNA_18 (.DIODE(_06763_));
 diode_2 ANTENNA_19 (.DIODE(_06763_));
 diode_2 ANTENNA_20 (.DIODE(_07098_));
 diode_2 ANTENNA_21 (.DIODE(_07113_));
 diode_2 ANTENNA_22 (.DIODE(_07852_));
 diode_2 ANTENNA_23 (.DIODE(_07852_));
 diode_2 ANTENNA_24 (.DIODE(_08527_));
 diode_2 ANTENNA_25 (.DIODE(_10095_));
 diode_2 ANTENNA_26 (.DIODE(_10417_));
 diode_2 ANTENNA_27 (.DIODE(_10814_));
 diode_2 ANTENNA_28 (.DIODE(_10830_));
 diode_2 ANTENNA_29 (.DIODE(_10830_));
 diode_2 ANTENNA_30 (.DIODE(_10840_));
 diode_2 ANTENNA_31 (.DIODE(_11110_));
 diode_2 ANTENNA_32 (.DIODE(clk_i));
 diode_2 ANTENNA_33 (.DIODE(\digitop_pav2.access_inst.access_check0.fg_i[0] ));
 diode_2 ANTENNA_34 (.DIODE(\digitop_pav2.access_inst.access_check0.fg_i[4] ));
 diode_2 ANTENNA_35 (.DIODE(\digitop_pav2.access_inst.access_check0.fg_i[8] ));
 diode_2 ANTENNA_36 (.DIODE(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[12] ));
 diode_2 ANTENNA_37 (.DIODE(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[12] ));
 diode_2 ANTENNA_38 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ));
 diode_2 ANTENNA_39 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state0_r[2] ));
 diode_2 ANTENNA_40 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ));
 diode_2 ANTENNA_41 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state1_r[11] ));
 diode_2 ANTENNA_42 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state1_r[2] ));
 diode_2 ANTENNA_43 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ));
 diode_2 ANTENNA_44 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ));
 diode_2 ANTENNA_45 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ));
 diode_2 ANTENNA_46 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state1_r[7] ));
 diode_2 ANTENNA_47 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state4_r[0] ));
 diode_2 ANTENNA_48 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state4_r[10] ));
 diode_2 ANTENNA_49 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state4_r[7] ));
 diode_2 ANTENNA_50 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state5_r[10] ));
 diode_2 ANTENNA_51 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state5_r[7] ));
 diode_2 ANTENNA_52 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state6_r[10] ));
 diode_2 ANTENNA_53 (.DIODE(\digitop_pav2.boot_inst.r_boot_ff ));
 diode_2 ANTENNA_54 (.DIODE(\digitop_pav2.func_clk ));
 diode_2 ANTENNA_55 (.DIODE(\digitop_pav2.func_clk ));
 diode_2 ANTENNA_56 (.DIODE(\digitop_pav2.func_rnclk_en ));
 diode_2 ANTENNA_57 (.DIODE(\digitop_pav2.invent_inst.invent_qqqr_pav2.sl_i ));
 diode_2 ANTENNA_58 (.DIODE(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[15] ));
 diode_2 ANTENNA_59 (.DIODE(\digitop_pav2.testctrl_pav2.inst_mbform.inst_form.int_rdata_i[15] ));
 diode_2 ANTENNA_60 (.DIODE(rnclk_i));
 diode_2 ANTENNA_61 (.DIODE(rnclk_i));
 diode_2 ANTENNA_62 (.DIODE(rnclk_i));
 diode_2 ANTENNA_63 (.DIODE(rnclk_i));
 diode_2 ANTENNA_64 (.DIODE(rr_data_i[20]));
 diode_2 ANTENNA_65 (.DIODE(rr_data_i[55]));
 diode_2 ANTENNA_66 (.DIODE(rr_data_i[63]));
 diode_2 ANTENNA_67 (.DIODE(\vmem_after_buf[111] ));
 diode_2 ANTENNA_68 (.DIODE(net13));
 diode_2 ANTENNA_69 (.DIODE(net16));
 diode_2 ANTENNA_70 (.DIODE(net21));
 diode_2 ANTENNA_71 (.DIODE(net21));
 diode_2 ANTENNA_72 (.DIODE(net22));
 diode_2 ANTENNA_73 (.DIODE(net25));
 diode_2 ANTENNA_74 (.DIODE(net67));
 diode_2 ANTENNA_75 (.DIODE(net67));
 diode_2 ANTENNA_76 (.DIODE(net84));
 diode_2 ANTENNA_77 (.DIODE(net84));
 diode_2 ANTENNA_78 (.DIODE(net84));
 diode_2 ANTENNA_79 (.DIODE(net84));
 diode_2 ANTENNA_80 (.DIODE(net84));
 diode_2 ANTENNA_81 (.DIODE(net84));
 diode_2 ANTENNA_82 (.DIODE(net84));
 diode_2 ANTENNA_83 (.DIODE(net84));
 diode_2 ANTENNA_84 (.DIODE(net84));
 diode_2 ANTENNA_85 (.DIODE(net84));
 diode_2 ANTENNA_86 (.DIODE(net85));
 diode_2 ANTENNA_87 (.DIODE(net85));
 diode_2 ANTENNA_88 (.DIODE(net85));
 diode_2 ANTENNA_89 (.DIODE(net85));
 diode_2 ANTENNA_90 (.DIODE(net85));
 diode_2 ANTENNA_91 (.DIODE(net85));
 diode_2 ANTENNA_92 (.DIODE(net85));
 diode_2 ANTENNA_93 (.DIODE(net85));
 diode_2 ANTENNA_94 (.DIODE(net85));
 diode_2 ANTENNA_95 (.DIODE(net85));
 diode_2 ANTENNA_96 (.DIODE(net86));
 diode_2 ANTENNA_97 (.DIODE(net87));
 diode_2 ANTENNA_98 (.DIODE(net87));
 diode_2 ANTENNA_99 (.DIODE(net87));
 diode_2 ANTENNA_100 (.DIODE(net87));
 diode_2 ANTENNA_101 (.DIODE(net87));
 diode_2 ANTENNA_102 (.DIODE(net87));
 diode_2 ANTENNA_103 (.DIODE(net89));
 diode_2 ANTENNA_104 (.DIODE(net95));
 diode_2 ANTENNA_105 (.DIODE(net95));
 diode_2 ANTENNA_106 (.DIODE(net103));
 diode_2 ANTENNA_107 (.DIODE(net103));
 diode_2 ANTENNA_108 (.DIODE(net105));
 diode_2 ANTENNA_109 (.DIODE(net301));
 diode_2 ANTENNA_110 (.DIODE(net308));
 diode_2 ANTENNA_111 (.DIODE(net308));
 diode_2 ANTENNA_112 (.DIODE(net313));
 diode_2 ANTENNA_113 (.DIODE(net313));
 diode_2 ANTENNA_114 (.DIODE(net313));
 diode_2 ANTENNA_115 (.DIODE(net313));
 diode_2 ANTENNA_116 (.DIODE(net313));
 diode_2 ANTENNA_117 (.DIODE(net313));
 diode_2 ANTENNA_118 (.DIODE(net313));
 diode_2 ANTENNA_119 (.DIODE(net313));
 diode_2 ANTENNA_120 (.DIODE(net313));
 diode_2 ANTENNA_121 (.DIODE(net313));
 diode_2 ANTENNA_122 (.DIODE(net314));
 diode_2 ANTENNA_123 (.DIODE(net314));
 diode_2 ANTENNA_124 (.DIODE(net314));
 diode_2 ANTENNA_125 (.DIODE(net412));
 diode_2 ANTENNA_126 (.DIODE(net675));
 diode_2 ANTENNA_127 (.DIODE(net675));
 diode_2 ANTENNA_128 (.DIODE(net729));
 diode_2 ANTENNA_129 (.DIODE(net905));
 diode_2 ANTENNA_130 (.DIODE(net911));
 diode_2 ANTENNA_131 (.DIODE(net955));
 diode_2 ANTENNA_132 (.DIODE(net1030));
 diode_2 ANTENNA_133 (.DIODE(net1086));
 diode_2 ANTENNA_134 (.DIODE(net1086));
 diode_2 ANTENNA_135 (.DIODE(net1086));
 diode_2 ANTENNA_136 (.DIODE(net1093));
 diode_2 ANTENNA_137 (.DIODE(net1095));
 diode_2 ANTENNA_138 (.DIODE(net1101));
 diode_2 ANTENNA_139 (.DIODE(net1105));
 diode_2 ANTENNA_140 (.DIODE(net1117));
 diode_2 ANTENNA_141 (.DIODE(net1119));
 diode_2 ANTENNA_142 (.DIODE(net1122));
 diode_2 ANTENNA_143 (.DIODE(net1123));
 diode_2 ANTENNA_144 (.DIODE(net1126));
 diode_2 ANTENNA_145 (.DIODE(net1133));
 diode_2 ANTENNA_146 (.DIODE(net1135));
 diode_2 ANTENNA_147 (.DIODE(net1135));
 diode_2 ANTENNA_148 (.DIODE(net1305));
 diode_2 ANTENNA_149 (.DIODE(net1322));
 diode_2 ANTENNA_150 (.DIODE(net1322));
 diode_2 ANTENNA_151 (.DIODE(net1457));
 diode_2 ANTENNA_152 (.DIODE(net1457));
 diode_2 ANTENNA_153 (.DIODE(net1503));
 diode_2 ANTENNA_154 (.DIODE(net1503));
 diode_2 ANTENNA_155 (.DIODE(net1503));
 diode_2 ANTENNA_156 (.DIODE(net1640));
 diode_2 ANTENNA_157 (.DIODE(net1640));
 diode_2 ANTENNA_158 (.DIODE(net1640));
 diode_2 ANTENNA_159 (.DIODE(net1640));
 diode_2 ANTENNA_160 (.DIODE(net1746));
 diode_2 ANTENNA_161 (.DIODE(_03308_));
 diode_2 ANTENNA_162 (.DIODE(_03701_));
 diode_2 ANTENNA_163 (.DIODE(_03759_));
 diode_2 ANTENNA_164 (.DIODE(_03760_));
 diode_2 ANTENNA_165 (.DIODE(_03760_));
 diode_2 ANTENNA_166 (.DIODE(_05622_));
 diode_2 ANTENNA_167 (.DIODE(_05788_));
 diode_2 ANTENNA_168 (.DIODE(_07061_));
 diode_2 ANTENNA_169 (.DIODE(_08928_));
 diode_2 ANTENNA_170 (.DIODE(_09537_));
 diode_2 ANTENNA_171 (.DIODE(\digitop_pav2.access_inst.access_check0.fg_i[2] ));
 diode_2 ANTENNA_172 (.DIODE(\digitop_pav2.access_inst.access_check0.permalock_tid_i ));
 diode_2 ANTENNA_173 (.DIODE(\digitop_pav2.access_inst.access_proc0.rd_dt_from_nvm_i[3] ));
 diode_2 ANTENNA_174 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state0_r[7] ));
 diode_2 ANTENNA_175 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state2_r[10] ));
 diode_2 ANTENNA_176 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state2_r[14] ));
 diode_2 ANTENNA_177 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state3_r[12] ));
 diode_2 ANTENNA_178 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state3_r[12] ));
 diode_2 ANTENNA_179 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state5_r[10] ));
 diode_2 ANTENNA_180 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state5_r[14] ));
 diode_2 ANTENNA_181 (.DIODE(\digitop_pav2.boot_inst.r_boot_ff ));
 diode_2 ANTENNA_182 (.DIODE(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ));
 diode_2 ANTENNA_183 (.DIODE(\digitop_pav2.invent_inst.invent_qqqr_pav2.s3_i ));
 diode_2 ANTENNA_184 (.DIODE(\digitop_pav2.memctrl_inst.addr_to_reram[3] ));
 diode_2 ANTENNA_185 (.DIODE(\digitop_pav2.proc_ctrl_inst.cmdfsm.n_rn_rst_b ));
 diode_2 ANTENNA_186 (.DIODE(\digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_i ));
 diode_2 ANTENNA_187 (.DIODE(\digitop_pav2.sync_inst.inst_clkx.inst_irreg.demod_i ));
 diode_2 ANTENNA_188 (.DIODE(rr_data_i[46]));
 diode_2 ANTENNA_189 (.DIODE(rr_data_i[47]));
 diode_2 ANTENNA_190 (.DIODE(\stadly_mpw03_erase_rise_9.Y ));
 diode_2 ANTENNA_191 (.DIODE(\vmem[383] ));
 diode_2 ANTENNA_192 (.DIODE(net10));
 diode_2 ANTENNA_193 (.DIODE(net26));
 diode_2 ANTENNA_194 (.DIODE(net34));
 diode_2 ANTENNA_195 (.DIODE(net53));
 diode_2 ANTENNA_196 (.DIODE(net68));
 diode_2 ANTENNA_197 (.DIODE(net159));
 diode_2 ANTENNA_198 (.DIODE(net309));
 diode_2 ANTENNA_199 (.DIODE(net309));
 diode_2 ANTENNA_200 (.DIODE(net459));
 diode_2 ANTENNA_201 (.DIODE(net470));
 diode_2 ANTENNA_202 (.DIODE(net648));
 diode_2 ANTENNA_203 (.DIODE(net648));
 diode_2 ANTENNA_204 (.DIODE(net648));
 diode_2 ANTENNA_205 (.DIODE(net648));
 diode_2 ANTENNA_206 (.DIODE(net800));
 diode_2 ANTENNA_207 (.DIODE(net1089));
 diode_2 ANTENNA_208 (.DIODE(net1089));
 diode_2 ANTENNA_209 (.DIODE(net1094));
 diode_2 ANTENNA_210 (.DIODE(net1123));
 diode_2 ANTENNA_211 (.DIODE(net1127));
 diode_2 ANTENNA_212 (.DIODE(net1483));
 diode_2 ANTENNA_213 (.DIODE(_06095_));
 diode_2 ANTENNA_214 (.DIODE(\digitop_pav2.aes128_inst.aes128_regs.state1_r[14] ));
 diode_2 ANTENNA_215 (.DIODE(rr_data_i[13]));
 diode_2 ANTENNA_216 (.DIODE(\vmem[11] ));
 diode_2 ANTENNA_217 (.DIODE(\vmem[63] ));
 diode_2 ANTENNA_218 (.DIODE(\vmem[95] ));
 diode_2 ANTENNA_219 (.DIODE(\vmem_after_buf[138] ));
 diode_2 ANTENNA_220 (.DIODE(\vmem_after_buf[90] ));
 diode_2 ANTENNA_221 (.DIODE(net723));
 diode_2 ANTENNA_222 (.DIODE(net769));
 diode_2 ANTENNA_223 (.DIODE(net1123));
 diode_2 ANTENNA_224 (.DIODE(net1324));
 decap_12 FILLER_0_9 ();
 fill_4 FILLER_0_21 ();
 fill_2 FILLER_0_25 ();
 fill_1 FILLER_0_27 ();
 fill_2 FILLER_0_32 ();
 fill_1 FILLER_0_34 ();
 fill_4 FILLER_0_39 ();
 fill_1 FILLER_0_43 ();
 fill_2 FILLER_0_50 ();
 fill_2 FILLER_0_65 ();
 fill_2 FILLER_0_95 ();
 fill_1 FILLER_0_106 ();
 fill_1 FILLER_0_111 ();
 fill_2 FILLER_0_113 ();
 fill_1 FILLER_0_115 ();
 fill_2 FILLER_0_123 ();
 fill_4 FILLER_0_128 ();
 fill_1 FILLER_0_132 ();
 fill_1 FILLER_0_139 ();
 fill_2 FILLER_0_141 ();
 fill_4 FILLER_0_155 ();
 fill_2 FILLER_0_159 ();
 fill_2 FILLER_0_165 ();
 fill_1 FILLER_0_167 ();
 fill_1 FILLER_0_169 ();
 fill_2 FILLER_0_174 ();
 fill_1 FILLER_0_176 ();
 fill_4 FILLER_0_183 ();
 fill_1 FILLER_0_187 ();
 fill_4 FILLER_0_192 ();
 fill_4 FILLER_0_201 ();
 fill_1 FILLER_0_205 ();
 fill_4 FILLER_0_210 ();
 fill_1 FILLER_0_214 ();
 fill_1 FILLER_0_219 ();
 fill_1 FILLER_0_247 ();
 fill_1 FILLER_0_253 ();
 fill_1 FILLER_0_270 ();
 fill_1 FILLER_0_279 ();
 fill_1 FILLER_0_281 ();
 fill_2 FILLER_0_290 ();
 fill_1 FILLER_0_318 ();
 fill_1 FILLER_0_355 ();
 fill_1 FILLER_0_365 ();
 fill_2 FILLER_0_474 ();
 fill_1 FILLER_0_497 ();
 fill_1 FILLER_0_559 ();
 fill_1 FILLER_0_587 ();
 fill_1 FILLER_0_595 ();
 fill_1 FILLER_0_623 ();
 fill_1 FILLER_0_633 ();
 fill_2 FILLER_0_698 ();
 fill_1 FILLER_0_727 ();
 fill_1 FILLER_0_729 ();
 fill_1 FILLER_0_785 ();
 fill_2 FILLER_0_810 ();
 fill_1 FILLER_0_833 ();
 fill_1 FILLER_0_863 ();
 fill_1 FILLER_0_886 ();
 fill_1 FILLER_0_903 ();
 fill_2 FILLER_0_953 ();
 fill_1 FILLER_0_979 ();
 fill_1 FILLER_0_1037 ();
 decap_12 FILLER_1_3 ();
 decap_12 FILLER_1_15 ();
 decap_12 FILLER_1_27 ();
 decap_12 FILLER_1_39 ();
 fill_4 FILLER_1_51 ();
 fill_1 FILLER_1_55 ();
 fill_2 FILLER_1_57 ();
 fill_2 FILLER_1_83 ();
 fill_1 FILLER_1_85 ();
 fill_1 FILLER_1_108 ();
 fill_2 FILLER_1_129 ();
 fill_2 FILLER_1_147 ();
 fill_2 FILLER_1_158 ();
 fill_4 FILLER_1_163 ();
 fill_1 FILLER_1_167 ();
 fill_4 FILLER_1_169 ();
 fill_1 FILLER_1_173 ();
 fill_4 FILLER_1_187 ();
 fill_1 FILLER_1_191 ();
 decap_12 FILLER_1_198 ();
 decap_12 FILLER_1_210 ();
 fill_2 FILLER_1_222 ();
 fill_4 FILLER_1_225 ();
 fill_1 FILLER_1_263 ();
 fill_1 FILLER_1_281 ();
 fill_1 FILLER_1_302 ();
 fill_2 FILLER_1_316 ();
 fill_2 FILLER_1_329 ();
 fill_1 FILLER_1_337 ();
 fill_1 FILLER_1_447 ();
 fill_2 FILLER_1_549 ();
 fill_2 FILLER_1_570 ();
 fill_4 FILLER_1_592 ();
 fill_2 FILLER_1_596 ();
 fill_1 FILLER_1_598 ();
 fill_2 FILLER_1_614 ();
 fill_2 FILLER_1_670 ();
 fill_1 FILLER_1_751 ();
 fill_1 FILLER_1_845 ();
 fill_1 FILLER_1_895 ();
 fill_1 FILLER_1_923 ();
 fill_2 FILLER_1_950 ();
 fill_1 FILLER_1_1029 ();
 decap_12 FILLER_2_3 ();
 decap_12 FILLER_2_15 ();
 fill_1 FILLER_2_27 ();
 decap_12 FILLER_2_29 ();
 fill_1 FILLER_2_41 ();
 fill_1 FILLER_2_62 ();
 fill_1 FILLER_2_83 ();
 fill_4 FILLER_2_85 ();
 fill_2 FILLER_2_89 ();
 fill_4 FILLER_2_100 ();
 fill_2 FILLER_2_104 ();
 decap_12 FILLER_2_109 ();
 fill_2 FILLER_2_121 ();
 decap_12 FILLER_2_126 ();
 fill_2 FILLER_2_138 ();
 fill_4 FILLER_2_141 ();
 fill_2 FILLER_2_145 ();
 decap_12 FILLER_2_152 ();
 fill_4 FILLER_2_164 ();
 fill_1 FILLER_2_168 ();
 fill_8 FILLER_2_172 ();
 fill_8 FILLER_2_188 ();
 decap_12 FILLER_2_197 ();
 decap_12 FILLER_2_209 ();
 fill_8 FILLER_2_221 ();
 fill_2 FILLER_2_229 ();
 fill_1 FILLER_2_231 ();
 fill_2 FILLER_2_235 ();
 fill_1 FILLER_2_237 ();
 fill_2 FILLER_2_267 ();
 fill_2 FILLER_2_273 ();
 fill_2 FILLER_2_290 ();
 fill_1 FILLER_2_307 ();
 fill_2 FILLER_2_309 ();
 fill_1 FILLER_2_322 ();
 fill_2 FILLER_2_365 ();
 fill_1 FILLER_2_376 ();
 fill_2 FILLER_2_506 ();
 fill_1 FILLER_2_533 ();
 fill_1 FILLER_2_643 ();
 fill_1 FILLER_2_645 ();
 fill_2 FILLER_2_710 ();
 fill_1 FILLER_2_749 ();
 fill_1 FILLER_2_793 ();
 fill_2 FILLER_2_866 ();
 fill_1 FILLER_2_882 ();
 fill_1 FILLER_2_969 ();
 fill_1 FILLER_2_979 ();
 fill_1 FILLER_2_1020 ();
 fill_1 FILLER_2_1037 ();
 decap_12 FILLER_3_3 ();
 decap_12 FILLER_3_15 ();
 decap_12 FILLER_3_27 ();
 decap_12 FILLER_3_39 ();
 fill_4 FILLER_3_51 ();
 fill_1 FILLER_3_55 ();
 decap_12 FILLER_3_57 ();
 fill_8 FILLER_3_69 ();
 fill_2 FILLER_3_77 ();
 fill_1 FILLER_3_79 ();
 fill_4 FILLER_3_85 ();
 fill_1 FILLER_3_89 ();
 decap_12 FILLER_3_95 ();
 fill_4 FILLER_3_107 ();
 fill_1 FILLER_3_111 ();
 fill_8 FILLER_3_113 ();
 fill_8 FILLER_3_126 ();
 fill_2 FILLER_3_148 ();
 fill_1 FILLER_3_150 ();
 fill_4 FILLER_3_154 ();
 fill_2 FILLER_3_158 ();
 decap_12 FILLER_3_177 ();
 fill_1 FILLER_3_189 ();
 decap_12 FILLER_3_210 ();
 fill_2 FILLER_3_222 ();
 fill_2 FILLER_3_225 ();
 fill_1 FILLER_3_227 ();
 fill_4 FILLER_3_237 ();
 fill_2 FILLER_3_278 ();
 fill_2 FILLER_3_300 ();
 fill_1 FILLER_3_320 ();
 fill_2 FILLER_3_334 ();
 fill_2 FILLER_3_337 ();
 fill_1 FILLER_3_384 ();
 fill_2 FILLER_3_505 ();
 fill_2 FILLER_3_621 ();
 fill_1 FILLER_3_671 ();
 fill_1 FILLER_3_673 ();
 fill_2 FILLER_3_710 ();
 fill_1 FILLER_3_721 ();
 fill_2 FILLER_3_738 ();
 fill_2 FILLER_3_809 ();
 fill_2 FILLER_3_829 ();
 fill_1 FILLER_3_895 ();
 fill_2 FILLER_3_930 ();
 fill_1 FILLER_3_956 ();
 fill_1 FILLER_3_1016 ();
 fill_1 FILLER_3_1037 ();
 decap_12 FILLER_4_3 ();
 decap_12 FILLER_4_15 ();
 fill_1 FILLER_4_27 ();
 decap_12 FILLER_4_29 ();
 decap_12 FILLER_4_41 ();
 fill_4 FILLER_4_53 ();
 fill_2 FILLER_4_57 ();
 fill_1 FILLER_4_59 ();
 fill_4 FILLER_4_80 ();
 fill_2 FILLER_4_90 ();
 fill_2 FILLER_4_100 ();
 fill_4 FILLER_4_115 ();
 fill_1 FILLER_4_119 ();
 fill_2 FILLER_4_148 ();
 fill_1 FILLER_4_150 ();
 decap_12 FILLER_4_161 ();
 fill_1 FILLER_4_173 ();
 fill_4 FILLER_4_190 ();
 fill_2 FILLER_4_194 ();
 fill_4 FILLER_4_197 ();
 fill_4 FILLER_4_211 ();
 fill_4 FILLER_4_232 ();
 fill_2 FILLER_4_236 ();
 fill_1 FILLER_4_251 ();
 fill_1 FILLER_4_260 ();
 fill_2 FILLER_4_267 ();
 fill_1 FILLER_4_269 ();
 fill_1 FILLER_4_281 ();
 fill_2 FILLER_4_306 ();
 fill_2 FILLER_4_309 ();
 fill_1 FILLER_4_335 ();
 fill_2 FILLER_4_347 ();
 fill_1 FILLER_4_365 ();
 fill_1 FILLER_4_382 ();
 fill_4 FILLER_4_397 ();
 fill_1 FILLER_4_401 ();
 fill_1 FILLER_4_433 ();
 fill_1 FILLER_4_521 ();
 fill_2 FILLER_4_533 ();
 fill_1 FILLER_4_587 ();
 fill_2 FILLER_4_633 ();
 fill_2 FILLER_4_645 ();
 fill_2 FILLER_4_676 ();
 fill_2 FILLER_4_707 ();
 fill_1 FILLER_4_709 ();
 fill_2 FILLER_4_866 ();
 fill_1 FILLER_4_889 ();
 fill_2 FILLER_4_904 ();
 fill_1 FILLER_4_934 ();
 fill_2 FILLER_4_1001 ();
 fill_2 FILLER_4_1015 ();
 fill_1 FILLER_4_1035 ();
 fill_1 FILLER_4_1037 ();
 decap_12 FILLER_5_3 ();
 fill_4 FILLER_5_15 ();
 decap_12 FILLER_5_40 ();
 fill_4 FILLER_5_52 ();
 decap_12 FILLER_5_57 ();
 decap_12 FILLER_5_69 ();
 fill_1 FILLER_5_81 ();
 decap_12 FILLER_5_87 ();
 decap_12 FILLER_5_99 ();
 fill_1 FILLER_5_111 ();
 fill_4 FILLER_5_113 ();
 fill_1 FILLER_5_117 ();
 fill_4 FILLER_5_124 ();
 fill_1 FILLER_5_128 ();
 decap_12 FILLER_5_148 ();
 fill_4 FILLER_5_160 ();
 fill_1 FILLER_5_164 ();
 fill_8 FILLER_5_177 ();
 fill_2 FILLER_5_185 ();
 fill_2 FILLER_5_194 ();
 decap_12 FILLER_5_199 ();
 decap_12 FILLER_5_211 ();
 fill_1 FILLER_5_223 ();
 decap_12 FILLER_5_225 ();
 fill_8 FILLER_5_237 ();
 fill_1 FILLER_5_245 ();
 fill_8 FILLER_5_249 ();
 fill_1 FILLER_5_257 ();
 decap_12 FILLER_5_268 ();
 fill_8 FILLER_5_281 ();
 fill_1 FILLER_5_292 ();
 fill_4 FILLER_5_296 ();
 fill_1 FILLER_5_300 ();
 fill_2 FILLER_5_312 ();
 fill_2 FILLER_5_322 ();
 fill_2 FILLER_5_342 ();
 fill_1 FILLER_5_393 ();
 fill_1 FILLER_5_443 ();
 fill_1 FILLER_5_492 ();
 fill_2 FILLER_5_502 ();
 fill_2 FILLER_5_505 ();
 fill_1 FILLER_5_516 ();
 fill_2 FILLER_5_549 ();
 fill_1 FILLER_5_567 ();
 fill_2 FILLER_5_588 ();
 fill_2 FILLER_5_605 ();
 fill_1 FILLER_5_617 ();
 fill_1 FILLER_5_633 ();
 fill_1 FILLER_5_671 ();
 fill_2 FILLER_5_682 ();
 fill_1 FILLER_5_721 ();
 fill_1 FILLER_5_729 ();
 fill_1 FILLER_5_744 ();
 fill_1 FILLER_5_783 ();
 fill_1 FILLER_5_839 ();
 fill_1 FILLER_5_845 ();
 fill_1 FILLER_5_876 ();
 fill_1 FILLER_5_895 ();
 fill_2 FILLER_5_900 ();
 fill_1 FILLER_5_926 ();
 fill_2 FILLER_5_950 ();
 fill_1 FILLER_5_962 ();
 fill_1 FILLER_5_993 ();
 fill_2 FILLER_5_1006 ();
 decap_12 FILLER_6_3 ();
 decap_12 FILLER_6_15 ();
 fill_1 FILLER_6_27 ();
 fill_4 FILLER_6_29 ();
 decap_12 FILLER_6_54 ();
 fill_8 FILLER_6_66 ();
 fill_2 FILLER_6_81 ();
 fill_1 FILLER_6_83 ();
 fill_2 FILLER_6_85 ();
 fill_4 FILLER_6_95 ();
 fill_4 FILLER_6_126 ();
 fill_1 FILLER_6_130 ();
 fill_1 FILLER_6_139 ();
 fill_4 FILLER_6_164 ();
 fill_1 FILLER_6_168 ();
 fill_4 FILLER_6_173 ();
 fill_2 FILLER_6_177 ();
 fill_1 FILLER_6_182 ();
 fill_1 FILLER_6_187 ();
 fill_1 FILLER_6_197 ();
 fill_8 FILLER_6_209 ();
 fill_1 FILLER_6_225 ();
 fill_4 FILLER_6_260 ();
 fill_4 FILLER_6_276 ();
 fill_2 FILLER_6_280 ();
 fill_4 FILLER_6_293 ();
 fill_2 FILLER_6_297 ();
 fill_4 FILLER_6_304 ();
 decap_12 FILLER_6_309 ();
 fill_4 FILLER_6_321 ();
 fill_2 FILLER_6_325 ();
 fill_2 FILLER_6_336 ();
 fill_2 FILLER_6_358 ();
 fill_2 FILLER_6_365 ();
 fill_1 FILLER_6_367 ();
 fill_4 FILLER_6_372 ();
 fill_1 FILLER_6_419 ();
 fill_2 FILLER_6_441 ();
 fill_1 FILLER_6_475 ();
 fill_2 FILLER_6_477 ();
 fill_2 FILLER_6_571 ();
 fill_1 FILLER_6_587 ();
 fill_2 FILLER_6_589 ();
 fill_2 FILLER_6_597 ();
 fill_1 FILLER_6_665 ();
 fill_1 FILLER_6_692 ();
 fill_1 FILLER_6_699 ();
 fill_1 FILLER_6_710 ();
 fill_1 FILLER_6_755 ();
 fill_1 FILLER_6_811 ();
 fill_2 FILLER_6_866 ();
 fill_2 FILLER_6_928 ();
 fill_2 FILLER_6_954 ();
 fill_1 FILLER_6_979 ();
 fill_2 FILLER_6_1019 ();
 fill_1 FILLER_6_1037 ();
 decap_12 FILLER_7_3 ();
 fill_8 FILLER_7_15 ();
 fill_1 FILLER_7_23 ();
 fill_1 FILLER_7_36 ();
 decap_12 FILLER_7_44 ();
 decap_12 FILLER_7_57 ();
 fill_1 FILLER_7_69 ();
 fill_8 FILLER_7_80 ();
 fill_1 FILLER_7_88 ();
 decap_12 FILLER_7_95 ();
 fill_4 FILLER_7_107 ();
 fill_1 FILLER_7_111 ();
 decap_12 FILLER_7_113 ();
 fill_4 FILLER_7_125 ();
 fill_1 FILLER_7_129 ();
 decap_12 FILLER_7_137 ();
 decap_12 FILLER_7_149 ();
 fill_1 FILLER_7_161 ();
 fill_2 FILLER_7_169 ();
 fill_1 FILLER_7_171 ();
 fill_4 FILLER_7_179 ();
 fill_2 FILLER_7_183 ();
 decap_12 FILLER_7_189 ();
 decap_12 FILLER_7_201 ();
 fill_4 FILLER_7_213 ();
 fill_2 FILLER_7_217 ();
 decap_12 FILLER_7_234 ();
 fill_4 FILLER_7_246 ();
 fill_1 FILLER_7_250 ();
 fill_2 FILLER_7_254 ();
 fill_8 FILLER_7_261 ();
 fill_2 FILLER_7_269 ();
 fill_2 FILLER_7_278 ();
 decap_12 FILLER_7_281 ();
 fill_1 FILLER_7_293 ();
 fill_1 FILLER_7_308 ();
 fill_8 FILLER_7_317 ();
 fill_2 FILLER_7_325 ();
 fill_1 FILLER_7_327 ();
 fill_1 FILLER_7_367 ();
 fill_1 FILLER_7_378 ();
 fill_1 FILLER_7_458 ();
 fill_1 FILLER_7_483 ();
 fill_1 FILLER_7_503 ();
 fill_2 FILLER_7_505 ();
 fill_2 FILLER_7_520 ();
 fill_1 FILLER_7_534 ();
 fill_2 FILLER_7_558 ();
 fill_2 FILLER_7_561 ();
 fill_2 FILLER_7_623 ();
 fill_1 FILLER_7_691 ();
 fill_1 FILLER_7_695 ();
 fill_1 FILLER_7_719 ();
 fill_2 FILLER_7_764 ();
 fill_2 FILLER_7_785 ();
 fill_2 FILLER_7_802 ();
 fill_1 FILLER_7_895 ();
 fill_2 FILLER_7_897 ();
 fill_1 FILLER_7_943 ();
 fill_2 FILLER_7_950 ();
 fill_1 FILLER_7_966 ();
 fill_1 FILLER_7_988 ();
 fill_1 FILLER_7_1007 ();
 fill_1 FILLER_7_1009 ();
 fill_2 FILLER_7_1036 ();
 decap_12 FILLER_8_7 ();
 fill_4 FILLER_8_19 ();
 fill_1 FILLER_8_23 ();
 fill_2 FILLER_8_38 ();
 fill_1 FILLER_8_40 ();
 fill_4 FILLER_8_68 ();
 fill_8 FILLER_8_75 ();
 fill_1 FILLER_8_83 ();
 fill_2 FILLER_8_96 ();
 fill_4 FILLER_8_114 ();
 fill_8 FILLER_8_121 ();
 fill_1 FILLER_8_129 ();
 fill_1 FILLER_8_139 ();
 fill_2 FILLER_8_141 ();
 fill_1 FILLER_8_143 ();
 decap_12 FILLER_8_151 ();
 fill_4 FILLER_8_166 ();
 fill_2 FILLER_8_170 ();
 fill_1 FILLER_8_172 ();
 decap_12 FILLER_8_176 ();
 fill_1 FILLER_8_188 ();
 fill_1 FILLER_8_195 ();
 decap_12 FILLER_8_200 ();
 fill_4 FILLER_8_212 ();
 fill_2 FILLER_8_216 ();
 fill_1 FILLER_8_218 ();
 fill_4 FILLER_8_230 ();
 fill_2 FILLER_8_250 ();
 fill_8 FILLER_8_261 ();
 fill_2 FILLER_8_269 ();
 fill_1 FILLER_8_271 ();
 decap_12 FILLER_8_285 ();
 fill_8 FILLER_8_297 ();
 fill_2 FILLER_8_305 ();
 fill_1 FILLER_8_307 ();
 fill_4 FILLER_8_309 ();
 decap_12 FILLER_8_322 ();
 fill_8 FILLER_8_334 ();
 fill_2 FILLER_8_345 ();
 fill_1 FILLER_8_347 ();
 fill_1 FILLER_8_357 ();
 fill_1 FILLER_8_380 ();
 fill_2 FILLER_8_402 ();
 fill_1 FILLER_8_419 ();
 fill_2 FILLER_8_421 ();
 fill_2 FILLER_8_444 ();
 fill_1 FILLER_8_475 ();
 fill_1 FILLER_8_500 ();
 fill_2 FILLER_8_530 ();
 fill_1 FILLER_8_533 ();
 fill_2 FILLER_8_589 ();
 fill_1 FILLER_8_631 ();
 fill_1 FILLER_8_645 ();
 fill_1 FILLER_8_678 ();
 fill_1 FILLER_8_682 ();
 fill_2 FILLER_8_692 ();
 fill_2 FILLER_8_701 ();
 fill_1 FILLER_8_715 ();
 fill_1 FILLER_8_787 ();
 fill_2 FILLER_8_866 ();
 fill_2 FILLER_8_925 ();
 fill_1 FILLER_8_979 ();
 fill_1 FILLER_8_990 ();
 fill_2 FILLER_8_1006 ();
 fill_1 FILLER_8_1035 ();
 fill_1 FILLER_8_1037 ();
 fill_2 FILLER_9_3 ();
 fill_1 FILLER_9_5 ();
 fill_1 FILLER_9_27 ();
 fill_1 FILLER_9_33 ();
 fill_2 FILLER_9_45 ();
 decap_12 FILLER_9_60 ();
 fill_4 FILLER_9_72 ();
 fill_2 FILLER_9_76 ();
 fill_1 FILLER_9_78 ();
 fill_2 FILLER_9_86 ();
 fill_1 FILLER_9_96 ();
 fill_4 FILLER_9_100 ();
 fill_2 FILLER_9_104 ();
 fill_1 FILLER_9_106 ();
 fill_2 FILLER_9_113 ();
 fill_1 FILLER_9_115 ();
 fill_2 FILLER_9_121 ();
 fill_1 FILLER_9_123 ();
 fill_4 FILLER_9_132 ();
 fill_1 FILLER_9_147 ();
 fill_2 FILLER_9_157 ();
 fill_1 FILLER_9_164 ();
 fill_2 FILLER_9_169 ();
 fill_1 FILLER_9_189 ();
 fill_2 FILLER_9_198 ();
 fill_4 FILLER_9_218 ();
 fill_2 FILLER_9_222 ();
 fill_1 FILLER_9_237 ();
 fill_4 FILLER_9_243 ();
 fill_2 FILLER_9_247 ();
 fill_1 FILLER_9_249 ();
 fill_1 FILLER_9_262 ();
 fill_1 FILLER_9_281 ();
 decap_12 FILLER_9_305 ();
 decap_12 FILLER_9_317 ();
 fill_4 FILLER_9_329 ();
 fill_2 FILLER_9_333 ();
 fill_1 FILLER_9_335 ();
 fill_1 FILLER_9_371 ();
 fill_2 FILLER_9_378 ();
 fill_1 FILLER_9_393 ();
 fill_1 FILLER_9_424 ();
 fill_2 FILLER_9_461 ();
 fill_1 FILLER_9_489 ();
 fill_2 FILLER_9_502 ();
 fill_1 FILLER_9_516 ();
 fill_2 FILLER_9_529 ();
 fill_2 FILLER_9_540 ();
 fill_1 FILLER_9_542 ();
 fill_2 FILLER_9_552 ();
 fill_2 FILLER_9_561 ();
 fill_1 FILLER_9_617 ();
 fill_1 FILLER_9_630 ();
 fill_1 FILLER_9_662 ();
 fill_1 FILLER_9_676 ();
 fill_2 FILLER_9_706 ();
 fill_1 FILLER_9_778 ();
 fill_1 FILLER_9_794 ();
 fill_1 FILLER_9_810 ();
 fill_1 FILLER_9_867 ();
 fill_1 FILLER_9_888 ();
 fill_1 FILLER_9_895 ();
 fill_2 FILLER_9_937 ();
 fill_1 FILLER_9_953 ();
 fill_2 FILLER_9_963 ();
 fill_1 FILLER_9_1015 ();
 fill_2 FILLER_9_1036 ();
 fill_4 FILLER_10_3 ();
 fill_4 FILLER_10_42 ();
 fill_8 FILLER_10_76 ();
 fill_4 FILLER_10_85 ();
 fill_2 FILLER_10_89 ();
 fill_1 FILLER_10_91 ();
 fill_4 FILLER_10_114 ();
 fill_2 FILLER_10_118 ();
 fill_1 FILLER_10_120 ();
 fill_4 FILLER_10_136 ();
 fill_4 FILLER_10_141 ();
 fill_1 FILLER_10_145 ();
 decap_12 FILLER_10_152 ();
 decap_12 FILLER_10_164 ();
 decap_12 FILLER_10_176 ();
 fill_4 FILLER_10_192 ();
 fill_8 FILLER_10_197 ();
 fill_1 FILLER_10_205 ();
 decap_12 FILLER_10_209 ();
 fill_2 FILLER_10_221 ();
 fill_1 FILLER_10_223 ();
 fill_4 FILLER_10_232 ();
 fill_2 FILLER_10_236 ();
 fill_4 FILLER_10_267 ();
 decap_12 FILLER_10_276 ();
 decap_12 FILLER_10_288 ();
 fill_1 FILLER_10_300 ();
 fill_4 FILLER_10_309 ();
 fill_2 FILLER_10_313 ();
 fill_1 FILLER_10_315 ();
 fill_4 FILLER_10_324 ();
 fill_1 FILLER_10_328 ();
 decap_12 FILLER_10_332 ();
 fill_4 FILLER_10_344 ();
 fill_2 FILLER_10_348 ();
 fill_1 FILLER_10_391 ();
 fill_2 FILLER_10_412 ();
 fill_4 FILLER_10_434 ();
 fill_1 FILLER_10_531 ();
 fill_2 FILLER_10_536 ();
 fill_1 FILLER_10_558 ();
 fill_2 FILLER_10_586 ();
 fill_1 FILLER_10_685 ();
 fill_2 FILLER_10_698 ();
 fill_2 FILLER_10_701 ();
 fill_1 FILLER_10_736 ();
 fill_1 FILLER_10_746 ();
 fill_1 FILLER_10_783 ();
 fill_1 FILLER_10_789 ();
 fill_2 FILLER_10_810 ();
 fill_1 FILLER_10_819 ();
 fill_2 FILLER_10_862 ();
 fill_1 FILLER_10_903 ();
 fill_2 FILLER_10_916 ();
 fill_2 FILLER_10_931 ();
 fill_1 FILLER_10_966 ();
 fill_1 FILLER_10_979 ();
 fill_1 FILLER_10_984 ();
 fill_1 FILLER_10_997 ();
 fill_2 FILLER_10_1030 ();
 fill_1 FILLER_10_1037 ();
 fill_8 FILLER_11_3 ();
 decap_12 FILLER_11_35 ();
 fill_1 FILLER_11_55 ();
 decap_12 FILLER_11_57 ();
 fill_2 FILLER_11_69 ();
 decap_12 FILLER_11_93 ();
 fill_4 FILLER_11_105 ();
 fill_1 FILLER_11_120 ();
 fill_2 FILLER_11_132 ();
 fill_2 FILLER_11_150 ();
 fill_2 FILLER_11_169 ();
 fill_2 FILLER_11_189 ();
 fill_4 FILLER_11_210 ();
 fill_4 FILLER_11_229 ();
 fill_2 FILLER_11_233 ();
 fill_1 FILLER_11_235 ();
 fill_4 FILLER_11_244 ();
 fill_1 FILLER_11_248 ();
 fill_2 FILLER_11_264 ();
 fill_1 FILLER_11_266 ();
 fill_2 FILLER_11_278 ();
 fill_2 FILLER_11_284 ();
 fill_4 FILLER_11_295 ();
 fill_4 FILLER_11_316 ();
 decap_12 FILLER_11_323 ();
 fill_1 FILLER_11_335 ();
 fill_2 FILLER_11_337 ();
 fill_4 FILLER_11_344 ();
 fill_1 FILLER_11_377 ();
 fill_1 FILLER_11_391 ();
 fill_1 FILLER_11_399 ();
 fill_1 FILLER_11_426 ();
 fill_2 FILLER_11_489 ();
 fill_1 FILLER_11_514 ();
 fill_8 FILLER_11_521 ();
 fill_2 FILLER_11_529 ();
 fill_1 FILLER_11_531 ();
 fill_1 FILLER_11_535 ();
 fill_1 FILLER_11_582 ();
 fill_4 FILLER_11_650 ();
 fill_2 FILLER_11_694 ();
 fill_1 FILLER_11_791 ();
 fill_1 FILLER_11_812 ();
 fill_1 FILLER_11_833 ();
 fill_2 FILLER_11_888 ();
 fill_2 FILLER_11_959 ();
 fill_1 FILLER_11_1007 ();
 fill_2 FILLER_11_1036 ();
 fill_4 FILLER_12_3 ();
 fill_2 FILLER_12_29 ();
 fill_2 FILLER_12_56 ();
 fill_2 FILLER_12_64 ();
 fill_1 FILLER_12_66 ();
 fill_1 FILLER_12_70 ();
 fill_8 FILLER_12_74 ();
 fill_2 FILLER_12_82 ();
 fill_4 FILLER_12_85 ();
 fill_1 FILLER_12_94 ();
 fill_4 FILLER_12_101 ();
 fill_1 FILLER_12_105 ();
 fill_4 FILLER_12_114 ();
 fill_1 FILLER_12_118 ();
 fill_1 FILLER_12_126 ();
 fill_1 FILLER_12_132 ();
 fill_2 FILLER_12_137 ();
 fill_1 FILLER_12_139 ();
 decap_12 FILLER_12_141 ();
 decap_12 FILLER_12_153 ();
 decap_12 FILLER_12_165 ();
 decap_12 FILLER_12_177 ();
 fill_4 FILLER_12_189 ();
 fill_2 FILLER_12_193 ();
 fill_1 FILLER_12_195 ();
 fill_2 FILLER_12_197 ();
 fill_1 FILLER_12_199 ();
 fill_8 FILLER_12_211 ();
 fill_1 FILLER_12_223 ();
 decap_12 FILLER_12_231 ();
 fill_8 FILLER_12_243 ();
 fill_1 FILLER_12_251 ();
 fill_4 FILLER_12_253 ();
 fill_1 FILLER_12_257 ();
 fill_8 FILLER_12_283 ();
 fill_4 FILLER_12_294 ();
 fill_2 FILLER_12_298 ();
 fill_1 FILLER_12_300 ();
 decap_12 FILLER_12_309 ();
 fill_4 FILLER_12_321 ();
 fill_2 FILLER_12_325 ();
 fill_1 FILLER_12_327 ();
 fill_2 FILLER_12_386 ();
 fill_2 FILLER_12_409 ();
 fill_2 FILLER_12_421 ();
 fill_1 FILLER_12_482 ();
 fill_2 FILLER_12_504 ();
 fill_2 FILLER_12_542 ();
 fill_1 FILLER_12_544 ();
 fill_2 FILLER_12_554 ();
 fill_1 FILLER_12_556 ();
 fill_2 FILLER_12_560 ();
 fill_1 FILLER_12_587 ();
 fill_1 FILLER_12_592 ();
 fill_2 FILLER_12_617 ();
 fill_4 FILLER_12_639 ();
 fill_1 FILLER_12_643 ();
 fill_2 FILLER_12_692 ();
 fill_1 FILLER_12_710 ();
 fill_1 FILLER_12_740 ();
 fill_2 FILLER_12_754 ();
 fill_1 FILLER_12_763 ();
 fill_2 FILLER_12_773 ();
 fill_2 FILLER_12_778 ();
 fill_1 FILLER_12_783 ();
 fill_2 FILLER_12_790 ();
 fill_4 FILLER_12_816 ();
 fill_2 FILLER_12_860 ();
 fill_1 FILLER_12_925 ();
 fill_2 FILLER_12_938 ();
 fill_2 FILLER_12_949 ();
 fill_1 FILLER_12_979 ();
 fill_1 FILLER_12_984 ();
 fill_2 FILLER_12_997 ();
 fill_1 FILLER_12_1008 ();
 fill_2 FILLER_12_1015 ();
 fill_1 FILLER_12_1029 ();
 fill_1 FILLER_12_1037 ();
 decap_12 FILLER_13_3 ();
 fill_2 FILLER_13_36 ();
 fill_4 FILLER_13_43 ();
 fill_2 FILLER_13_47 ();
 fill_2 FILLER_13_54 ();
 fill_4 FILLER_13_60 ();
 fill_1 FILLER_13_64 ();
 fill_8 FILLER_13_73 ();
 fill_1 FILLER_13_81 ();
 fill_2 FILLER_13_113 ();
 fill_1 FILLER_13_115 ();
 decap_12 FILLER_13_143 ();
 fill_4 FILLER_13_155 ();
 fill_2 FILLER_13_159 ();
 fill_1 FILLER_13_161 ();
 fill_2 FILLER_13_165 ();
 fill_1 FILLER_13_167 ();
 fill_2 FILLER_13_169 ();
 fill_4 FILLER_13_179 ();
 fill_2 FILLER_13_183 ();
 fill_4 FILLER_13_193 ();
 fill_2 FILLER_13_197 ();
 fill_1 FILLER_13_199 ();
 fill_4 FILLER_13_217 ();
 fill_2 FILLER_13_221 ();
 fill_1 FILLER_13_223 ();
 fill_1 FILLER_13_225 ();
 fill_4 FILLER_13_244 ();
 fill_2 FILLER_13_248 ();
 fill_2 FILLER_13_266 ();
 fill_4 FILLER_13_275 ();
 fill_1 FILLER_13_279 ();
 fill_4 FILLER_13_281 ();
 fill_2 FILLER_13_285 ();
 fill_1 FILLER_13_287 ();
 fill_8 FILLER_13_325 ();
 fill_2 FILLER_13_333 ();
 fill_1 FILLER_13_335 ();
 fill_8 FILLER_13_345 ();
 fill_1 FILLER_13_353 ();
 fill_1 FILLER_13_483 ();
 fill_1 FILLER_13_505 ();
 fill_2 FILLER_13_521 ();
 fill_2 FILLER_13_529 ();
 fill_1 FILLER_13_531 ();
 fill_4 FILLER_13_535 ();
 fill_1 FILLER_13_559 ();
 fill_2 FILLER_13_613 ();
 fill_1 FILLER_13_615 ();
 fill_2 FILLER_13_632 ();
 fill_1 FILLER_13_634 ();
 fill_1 FILLER_13_638 ();
 fill_2 FILLER_13_670 ();
 fill_1 FILLER_13_694 ();
 fill_2 FILLER_13_738 ();
 fill_2 FILLER_13_811 ();
 fill_2 FILLER_13_885 ();
 fill_1 FILLER_13_922 ();
 fill_1 FILLER_13_963 ();
 fill_1 FILLER_13_979 ();
 decap_12 FILLER_14_3 ();
 decap_12 FILLER_14_15 ();
 fill_1 FILLER_14_27 ();
 fill_1 FILLER_14_29 ();
 fill_1 FILLER_14_65 ();
 fill_4 FILLER_14_70 ();
 fill_1 FILLER_14_74 ();
 fill_2 FILLER_14_81 ();
 fill_1 FILLER_14_83 ();
 decap_12 FILLER_14_85 ();
 fill_2 FILLER_14_97 ();
 fill_1 FILLER_14_99 ();
 fill_4 FILLER_14_106 ();
 fill_2 FILLER_14_110 ();
 fill_1 FILLER_14_112 ();
 fill_4 FILLER_14_136 ();
 fill_1 FILLER_14_141 ();
 fill_2 FILLER_14_167 ();
 fill_1 FILLER_14_180 ();
 fill_2 FILLER_14_193 ();
 fill_1 FILLER_14_195 ();
 fill_4 FILLER_14_201 ();
 fill_2 FILLER_14_205 ();
 fill_4 FILLER_14_210 ();
 fill_1 FILLER_14_214 ();
 fill_2 FILLER_14_222 ();
 fill_2 FILLER_14_236 ();
 fill_1 FILLER_14_238 ();
 fill_4 FILLER_14_248 ();
 fill_4 FILLER_14_253 ();
 fill_2 FILLER_14_257 ();
 fill_1 FILLER_14_259 ();
 fill_4 FILLER_14_268 ();
 fill_1 FILLER_14_272 ();
 fill_1 FILLER_14_315 ();
 decap_12 FILLER_14_323 ();
 fill_1 FILLER_14_335 ();
 decap_12 FILLER_14_347 ();
 fill_4 FILLER_14_359 ();
 fill_1 FILLER_14_363 ();
 fill_4 FILLER_14_365 ();
 fill_1 FILLER_14_369 ();
 fill_1 FILLER_14_389 ();
 fill_1 FILLER_14_419 ();
 fill_2 FILLER_14_421 ();
 fill_1 FILLER_14_438 ();
 fill_2 FILLER_14_459 ();
 fill_1 FILLER_14_461 ();
 fill_2 FILLER_14_477 ();
 fill_2 FILLER_14_511 ();
 fill_1 FILLER_14_513 ();
 fill_2 FILLER_14_518 ();
 fill_4 FILLER_14_538 ();
 fill_2 FILLER_14_558 ();
 fill_1 FILLER_14_579 ();
 fill_2 FILLER_14_586 ();
 fill_1 FILLER_14_598 ();
 fill_4 FILLER_14_605 ();
 fill_1 FILLER_14_609 ();
 fill_4 FILLER_14_640 ();
 fill_1 FILLER_14_651 ();
 fill_2 FILLER_14_664 ();
 fill_1 FILLER_14_699 ();
 fill_2 FILLER_14_710 ();
 fill_2 FILLER_14_773 ();
 fill_2 FILLER_14_784 ();
 fill_1 FILLER_14_795 ();
 fill_1 FILLER_14_811 ();
 fill_1 FILLER_14_904 ();
 fill_2 FILLER_14_922 ();
 fill_2 FILLER_14_955 ();
 fill_2 FILLER_14_981 ();
 fill_1 FILLER_14_992 ();
 fill_2 FILLER_14_1024 ();
 fill_1 FILLER_14_1035 ();
 fill_1 FILLER_14_1037 ();
 decap_12 FILLER_15_3 ();
 fill_2 FILLER_15_15 ();
 fill_4 FILLER_15_51 ();
 fill_1 FILLER_15_55 ();
 decap_12 FILLER_15_57 ();
 fill_4 FILLER_15_69 ();
 fill_2 FILLER_15_73 ();
 fill_4 FILLER_15_82 ();
 fill_1 FILLER_15_86 ();
 fill_2 FILLER_15_109 ();
 fill_1 FILLER_15_111 ();
 fill_2 FILLER_15_143 ();
 fill_1 FILLER_15_145 ();
 fill_4 FILLER_15_161 ();
 fill_2 FILLER_15_165 ();
 fill_1 FILLER_15_167 ();
 fill_8 FILLER_15_169 ();
 fill_1 FILLER_15_177 ();
 fill_2 FILLER_15_193 ();
 fill_1 FILLER_15_206 ();
 fill_1 FILLER_15_223 ();
 fill_2 FILLER_15_263 ();
 fill_1 FILLER_15_265 ();
 fill_4 FILLER_15_275 ();
 fill_1 FILLER_15_279 ();
 fill_1 FILLER_15_289 ();
 fill_2 FILLER_15_298 ();
 fill_4 FILLER_15_317 ();
 fill_2 FILLER_15_321 ();
 fill_1 FILLER_15_327 ();
 fill_2 FILLER_15_333 ();
 fill_1 FILLER_15_335 ();
 fill_4 FILLER_15_337 ();
 decap_12 FILLER_15_344 ();
 fill_2 FILLER_15_356 ();
 fill_2 FILLER_15_378 ();
 fill_1 FILLER_15_380 ();
 fill_4 FILLER_15_386 ();
 fill_2 FILLER_15_390 ();
 fill_2 FILLER_15_393 ();
 fill_1 FILLER_15_395 ();
 fill_4 FILLER_15_399 ();
 fill_2 FILLER_15_403 ();
 fill_2 FILLER_15_429 ();
 fill_2 FILLER_15_434 ();
 fill_1 FILLER_15_436 ();
 fill_8 FILLER_15_440 ();
 fill_4 FILLER_15_455 ();
 fill_2 FILLER_15_459 ();
 fill_2 FILLER_15_481 ();
 fill_1 FILLER_15_505 ();
 fill_2 FILLER_15_535 ();
 fill_1 FILLER_15_552 ();
 fill_1 FILLER_15_556 ();
 fill_4 FILLER_15_599 ();
 fill_2 FILLER_15_603 ();
 fill_2 FILLER_15_614 ();
 fill_1 FILLER_15_656 ();
 fill_1 FILLER_15_671 ();
 fill_2 FILLER_15_726 ();
 fill_1 FILLER_15_794 ();
 fill_1 FILLER_15_839 ();
 fill_2 FILLER_15_894 ();
 fill_2 FILLER_15_897 ();
 fill_1 FILLER_15_951 ();
 fill_2 FILLER_15_989 ();
 fill_2 FILLER_15_1003 ();
 decap_12 FILLER_16_3 ();
 decap_12 FILLER_16_15 ();
 fill_1 FILLER_16_27 ();
 fill_2 FILLER_16_29 ();
 fill_1 FILLER_16_31 ();
 fill_8 FILLER_16_74 ();
 fill_2 FILLER_16_82 ();
 fill_8 FILLER_16_93 ();
 fill_4 FILLER_16_111 ();
 fill_2 FILLER_16_115 ();
 fill_8 FILLER_16_125 ();
 fill_2 FILLER_16_133 ();
 fill_1 FILLER_16_135 ();
 fill_2 FILLER_16_145 ();
 fill_1 FILLER_16_147 ();
 fill_4 FILLER_16_151 ();
 fill_1 FILLER_16_155 ();
 fill_1 FILLER_16_163 ();
 fill_1 FILLER_16_181 ();
 fill_2 FILLER_16_211 ();
 fill_1 FILLER_16_221 ();
 fill_2 FILLER_16_226 ();
 fill_1 FILLER_16_228 ();
 fill_1 FILLER_16_244 ();
 fill_2 FILLER_16_265 ();
 fill_1 FILLER_16_267 ();
 fill_4 FILLER_16_272 ();
 fill_2 FILLER_16_276 ();
 fill_8 FILLER_16_287 ();
 fill_1 FILLER_16_295 ();
 fill_4 FILLER_16_301 ();
 fill_2 FILLER_16_305 ();
 fill_1 FILLER_16_307 ();
 fill_2 FILLER_16_318 ();
 fill_4 FILLER_16_334 ();
 fill_1 FILLER_16_343 ();
 fill_4 FILLER_16_350 ();
 fill_2 FILLER_16_354 ();
 fill_1 FILLER_16_363 ();
 fill_8 FILLER_16_365 ();
 fill_2 FILLER_16_373 ();
 fill_1 FILLER_16_419 ();
 decap_12 FILLER_16_424 ();
 fill_2 FILLER_16_436 ();
 fill_4 FILLER_16_472 ();
 fill_2 FILLER_16_483 ();
 fill_2 FILLER_16_517 ();
 fill_1 FILLER_16_519 ();
 fill_2 FILLER_16_533 ();
 fill_1 FILLER_16_535 ();
 fill_2 FILLER_16_690 ();
 fill_1 FILLER_16_705 ();
 fill_4 FILLER_16_751 ();
 fill_1 FILLER_16_755 ();
 fill_1 FILLER_16_779 ();
 fill_1 FILLER_16_813 ();
 fill_2 FILLER_16_827 ();
 fill_2 FILLER_16_849 ();
 fill_1 FILLER_16_851 ();
 fill_1 FILLER_16_869 ();
 fill_1 FILLER_16_879 ();
 fill_1 FILLER_16_895 ();
 fill_2 FILLER_16_978 ();
 fill_1 FILLER_16_1037 ();
 decap_12 FILLER_17_3 ();
 fill_4 FILLER_17_15 ();
 fill_2 FILLER_17_19 ();
 fill_2 FILLER_17_50 ();
 fill_4 FILLER_17_83 ();
 fill_1 FILLER_17_87 ();
 fill_4 FILLER_17_106 ();
 fill_2 FILLER_17_110 ();
 fill_2 FILLER_17_121 ();
 fill_1 FILLER_17_123 ();
 decap_12 FILLER_17_130 ();
 fill_1 FILLER_17_142 ();
 fill_2 FILLER_17_150 ();
 fill_4 FILLER_17_169 ();
 fill_2 FILLER_17_173 ();
 fill_1 FILLER_17_175 ();
 fill_8 FILLER_17_182 ();
 fill_2 FILLER_17_190 ();
 fill_1 FILLER_17_192 ();
 fill_4 FILLER_17_206 ();
 fill_2 FILLER_17_210 ();
 fill_1 FILLER_17_212 ();
 fill_4 FILLER_17_220 ();
 fill_4 FILLER_17_254 ();
 fill_2 FILLER_17_266 ();
 fill_1 FILLER_17_268 ();
 fill_4 FILLER_17_289 ();
 fill_1 FILLER_17_293 ();
 fill_4 FILLER_17_302 ();
 fill_2 FILLER_17_306 ();
 fill_1 FILLER_17_308 ();
 fill_4 FILLER_17_320 ();
 fill_1 FILLER_17_324 ();
 fill_4 FILLER_17_330 ();
 fill_2 FILLER_17_334 ();
 fill_2 FILLER_17_337 ();
 fill_4 FILLER_17_342 ();
 fill_2 FILLER_17_346 ();
 fill_1 FILLER_17_378 ();
 fill_2 FILLER_17_382 ();
 fill_1 FILLER_17_418 ();
 fill_1 FILLER_17_447 ();
 fill_2 FILLER_17_449 ();
 fill_1 FILLER_17_451 ();
 fill_1 FILLER_17_468 ();
 fill_1 FILLER_17_505 ();
 fill_1 FILLER_17_550 ();
 fill_2 FILLER_17_579 ();
 fill_1 FILLER_17_604 ();
 fill_2 FILLER_17_611 ();
 fill_1 FILLER_17_631 ();
 fill_2 FILLER_17_655 ();
 fill_4 FILLER_17_665 ();
 fill_2 FILLER_17_669 ();
 fill_1 FILLER_17_671 ();
 fill_2 FILLER_17_673 ();
 fill_1 FILLER_17_675 ();
 fill_2 FILLER_17_755 ();
 fill_1 FILLER_17_783 ();
 fill_1 FILLER_17_796 ();
 fill_1 FILLER_17_839 ();
 fill_2 FILLER_17_844 ();
 fill_2 FILLER_17_866 ();
 fill_2 FILLER_17_874 ();
 fill_2 FILLER_17_913 ();
 fill_1 FILLER_17_935 ();
 fill_1 FILLER_17_942 ();
 fill_1 FILLER_17_996 ();
 fill_2 FILLER_17_1006 ();
 fill_2 FILLER_17_1036 ();
 decap_12 FILLER_18_3 ();
 fill_8 FILLER_18_15 ();
 fill_1 FILLER_18_23 ();
 fill_2 FILLER_18_44 ();
 fill_1 FILLER_18_46 ();
 fill_4 FILLER_18_67 ();
 fill_2 FILLER_18_71 ();
 fill_1 FILLER_18_73 ();
 fill_4 FILLER_18_77 ();
 fill_2 FILLER_18_81 ();
 fill_1 FILLER_18_83 ();
 fill_1 FILLER_18_85 ();
 decap_12 FILLER_18_90 ();
 decap_12 FILLER_18_102 ();
 fill_2 FILLER_18_114 ();
 fill_4 FILLER_18_125 ();
 fill_2 FILLER_18_129 ();
 fill_1 FILLER_18_131 ();
 fill_2 FILLER_18_138 ();
 fill_4 FILLER_18_141 ();
 fill_1 FILLER_18_145 ();
 fill_2 FILLER_18_149 ();
 decap_12 FILLER_18_154 ();
 fill_8 FILLER_18_166 ();
 fill_2 FILLER_18_174 ();
 fill_4 FILLER_18_183 ();
 fill_1 FILLER_18_187 ();
 fill_2 FILLER_18_197 ();
 fill_1 FILLER_18_210 ();
 fill_4 FILLER_18_219 ();
 fill_2 FILLER_18_238 ();
 fill_4 FILLER_18_261 ();
 fill_2 FILLER_18_265 ();
 fill_8 FILLER_18_274 ();
 fill_2 FILLER_18_282 ();
 fill_1 FILLER_18_284 ();
 decap_12 FILLER_18_288 ();
 fill_4 FILLER_18_303 ();
 fill_1 FILLER_18_307 ();
 fill_1 FILLER_18_322 ();
 fill_8 FILLER_18_328 ();
 fill_1 FILLER_18_336 ();
 fill_2 FILLER_18_347 ();
 fill_1 FILLER_18_349 ();
 fill_2 FILLER_18_362 ();
 fill_2 FILLER_18_412 ();
 fill_4 FILLER_18_421 ();
 fill_2 FILLER_18_425 ();
 fill_1 FILLER_18_427 ();
 fill_2 FILLER_18_437 ();
 fill_2 FILLER_18_451 ();
 fill_2 FILLER_18_464 ();
 fill_2 FILLER_18_474 ();
 fill_1 FILLER_18_533 ();
 fill_2 FILLER_18_553 ();
 fill_1 FILLER_18_555 ();
 fill_2 FILLER_18_589 ();
 fill_1 FILLER_18_615 ();
 fill_1 FILLER_18_645 ();
 fill_1 FILLER_18_662 ();
 fill_4 FILLER_18_666 ();
 fill_2 FILLER_18_670 ();
 fill_1 FILLER_18_672 ();
 fill_1 FILLER_18_680 ();
 fill_4 FILLER_18_688 ();
 fill_1 FILLER_18_692 ();
 fill_2 FILLER_18_707 ();
 fill_2 FILLER_18_741 ();
 fill_1 FILLER_18_811 ();
 fill_2 FILLER_18_849 ();
 fill_2 FILLER_18_857 ();
 fill_2 FILLER_18_931 ();
 fill_1 FILLER_18_979 ();
 fill_1 FILLER_18_1029 ();
 fill_1 FILLER_18_1037 ();
 fill_4 FILLER_19_3 ();
 fill_1 FILLER_19_7 ();
 fill_2 FILLER_19_54 ();
 fill_2 FILLER_19_57 ();
 fill_1 FILLER_19_59 ();
 decap_12 FILLER_19_71 ();
 fill_4 FILLER_19_83 ();
 fill_2 FILLER_19_87 ();
 fill_1 FILLER_19_89 ();
 fill_4 FILLER_19_99 ();
 fill_4 FILLER_19_108 ();
 fill_8 FILLER_19_113 ();
 fill_2 FILLER_19_121 ();
 fill_2 FILLER_19_130 ();
 fill_2 FILLER_19_156 ();
 fill_2 FILLER_19_162 ();
 fill_1 FILLER_19_164 ();
 fill_1 FILLER_19_176 ();
 fill_4 FILLER_19_182 ();
 fill_2 FILLER_19_186 ();
 decap_12 FILLER_19_194 ();
 fill_8 FILLER_19_206 ();
 fill_1 FILLER_19_214 ();
 fill_2 FILLER_19_221 ();
 fill_1 FILLER_19_223 ();
 fill_1 FILLER_19_230 ();
 decap_12 FILLER_19_234 ();
 fill_4 FILLER_19_246 ();
 fill_1 FILLER_19_250 ();
 fill_1 FILLER_19_262 ();
 fill_2 FILLER_19_266 ();
 fill_4 FILLER_19_273 ();
 fill_2 FILLER_19_277 ();
 fill_1 FILLER_19_279 ();
 fill_1 FILLER_19_281 ();
 decap_12 FILLER_19_318 ();
 fill_4 FILLER_19_330 ();
 fill_2 FILLER_19_334 ();
 fill_2 FILLER_19_345 ();
 fill_2 FILLER_19_368 ();
 fill_2 FILLER_19_390 ();
 fill_1 FILLER_19_447 ();
 fill_1 FILLER_19_470 ();
 fill_1 FILLER_19_485 ();
 fill_1 FILLER_19_489 ();
 fill_2 FILLER_19_499 ();
 fill_1 FILLER_19_525 ();
 fill_2 FILLER_19_561 ();
 fill_1 FILLER_19_563 ();
 fill_1 FILLER_19_626 ();
 fill_1 FILLER_19_673 ();
 fill_1 FILLER_19_694 ();
 fill_4 FILLER_19_701 ();
 fill_2 FILLER_19_705 ();
 fill_1 FILLER_19_720 ();
 fill_2 FILLER_19_732 ();
 fill_2 FILLER_19_763 ();
 fill_2 FILLER_19_807 ();
 fill_1 FILLER_19_818 ();
 fill_1 FILLER_19_920 ();
 fill_1 FILLER_19_951 ();
 fill_1 FILLER_19_988 ();
 fill_1 FILLER_19_1004 ();
 fill_2 FILLER_19_1009 ();
 decap_12 FILLER_20_3 ();
 fill_4 FILLER_20_15 ();
 fill_2 FILLER_20_19 ();
 fill_1 FILLER_20_21 ();
 fill_4 FILLER_20_29 ();
 fill_1 FILLER_20_39 ();
 fill_4 FILLER_20_45 ();
 fill_1 FILLER_20_49 ();
 fill_4 FILLER_20_56 ();
 fill_4 FILLER_20_80 ();
 fill_1 FILLER_20_92 ();
 fill_2 FILLER_20_99 ();
 fill_1 FILLER_20_101 ();
 fill_2 FILLER_20_116 ();
 fill_1 FILLER_20_118 ();
 decap_12 FILLER_20_126 ();
 fill_2 FILLER_20_138 ();
 decap_12 FILLER_20_141 ();
 decap_12 FILLER_20_158 ();
 fill_1 FILLER_20_170 ();
 fill_4 FILLER_20_179 ();
 fill_2 FILLER_20_183 ();
 fill_1 FILLER_20_195 ();
 fill_4 FILLER_20_197 ();
 fill_1 FILLER_20_201 ();
 fill_2 FILLER_20_212 ();
 fill_1 FILLER_20_214 ();
 fill_2 FILLER_20_233 ();
 fill_2 FILLER_20_249 ();
 fill_1 FILLER_20_251 ();
 fill_8 FILLER_20_265 ();
 fill_2 FILLER_20_273 ();
 fill_4 FILLER_20_279 ();
 fill_2 FILLER_20_296 ();
 fill_1 FILLER_20_298 ();
 fill_2 FILLER_20_306 ();
 fill_2 FILLER_20_315 ();
 fill_1 FILLER_20_336 ();
 fill_1 FILLER_20_343 ();
 fill_1 FILLER_20_365 ();
 decap_12 FILLER_20_396 ();
 fill_4 FILLER_20_408 ();
 fill_2 FILLER_20_412 ();
 fill_2 FILLER_20_418 ();
 fill_8 FILLER_20_421 ();
 fill_2 FILLER_20_429 ();
 fill_4 FILLER_20_434 ();
 fill_1 FILLER_20_438 ();
 fill_2 FILLER_20_465 ();
 fill_2 FILLER_20_542 ();
 fill_1 FILLER_20_544 ();
 fill_1 FILLER_20_554 ();
 fill_2 FILLER_20_651 ();
 fill_2 FILLER_20_671 ();
 fill_4 FILLER_20_693 ();
 fill_2 FILLER_20_697 ();
 fill_1 FILLER_20_699 ();
 decap_12 FILLER_20_721 ();
 fill_2 FILLER_20_746 ();
 fill_2 FILLER_20_754 ();
 fill_1 FILLER_20_792 ();
 fill_1 FILLER_20_867 ();
 fill_1 FILLER_20_882 ();
 fill_1 FILLER_20_889 ();
 fill_1 FILLER_20_945 ();
 fill_2 FILLER_20_978 ();
 fill_1 FILLER_20_1035 ();
 fill_1 FILLER_20_1037 ();
 fill_8 FILLER_21_3 ();
 fill_2 FILLER_21_11 ();
 fill_1 FILLER_21_18 ();
 fill_2 FILLER_21_22 ();
 fill_1 FILLER_21_24 ();
 fill_2 FILLER_21_30 ();
 fill_1 FILLER_21_32 ();
 fill_8 FILLER_21_38 ();
 fill_8 FILLER_21_57 ();
 fill_2 FILLER_21_65 ();
 fill_1 FILLER_21_67 ();
 decap_12 FILLER_21_71 ();
 fill_8 FILLER_21_83 ();
 fill_8 FILLER_21_104 ();
 fill_2 FILLER_21_113 ();
 fill_1 FILLER_21_115 ();
 fill_2 FILLER_21_128 ();
 fill_2 FILLER_21_147 ();
 fill_1 FILLER_21_169 ();
 fill_1 FILLER_21_173 ();
 fill_4 FILLER_21_186 ();
 decap_12 FILLER_21_198 ();
 fill_2 FILLER_21_210 ();
 fill_4 FILLER_21_219 ();
 fill_1 FILLER_21_223 ();
 fill_8 FILLER_21_225 ();
 fill_2 FILLER_21_233 ();
 fill_1 FILLER_21_238 ();
 fill_4 FILLER_21_242 ();
 fill_2 FILLER_21_246 ();
 fill_1 FILLER_21_248 ();
 fill_8 FILLER_21_255 ();
 fill_1 FILLER_21_263 ();
 fill_1 FILLER_21_270 ();
 fill_2 FILLER_21_277 ();
 fill_1 FILLER_21_279 ();
 fill_2 FILLER_21_281 ();
 fill_8 FILLER_21_290 ();
 fill_8 FILLER_21_301 ();
 fill_2 FILLER_21_309 ();
 fill_1 FILLER_21_311 ();
 decap_12 FILLER_21_319 ();
 fill_4 FILLER_21_331 ();
 fill_1 FILLER_21_335 ();
 decap_12 FILLER_21_337 ();
 fill_8 FILLER_21_349 ();
 fill_1 FILLER_21_377 ();
 fill_1 FILLER_21_385 ();
 fill_2 FILLER_21_389 ();
 fill_1 FILLER_21_391 ();
 fill_2 FILLER_21_413 ();
 fill_4 FILLER_21_443 ();
 fill_1 FILLER_21_447 ();
 fill_4 FILLER_21_449 ();
 fill_1 FILLER_21_453 ();
 fill_2 FILLER_21_487 ();
 fill_2 FILLER_21_502 ();
 fill_2 FILLER_21_505 ();
 fill_1 FILLER_21_516 ();
 fill_4 FILLER_21_529 ();
 fill_1 FILLER_21_559 ();
 fill_1 FILLER_21_623 ();
 fill_1 FILLER_21_640 ();
 fill_1 FILLER_21_671 ();
 fill_4 FILLER_21_681 ();
 fill_1 FILLER_21_685 ();
 fill_4 FILLER_21_723 ();
 fill_1 FILLER_21_727 ();
 fill_1 FILLER_21_736 ();
 fill_1 FILLER_21_754 ();
 fill_1 FILLER_21_818 ();
 fill_1 FILLER_21_839 ();
 fill_2 FILLER_21_850 ();
 fill_1 FILLER_21_957 ();
 fill_2 FILLER_21_987 ();
 fill_2 FILLER_21_1033 ();
 fill_4 FILLER_22_3 ();
 fill_2 FILLER_22_7 ();
 decap_12 FILLER_22_16 ();
 fill_4 FILLER_22_38 ();
 fill_1 FILLER_22_47 ();
 fill_8 FILLER_22_51 ();
 fill_1 FILLER_22_70 ();
 fill_8 FILLER_22_74 ();
 fill_2 FILLER_22_82 ();
 fill_4 FILLER_22_88 ();
 fill_2 FILLER_22_123 ();
 fill_8 FILLER_22_131 ();
 fill_1 FILLER_22_139 ();
 decap_12 FILLER_22_141 ();
 fill_4 FILLER_22_153 ();
 fill_2 FILLER_22_157 ();
 fill_8 FILLER_22_163 ();
 fill_2 FILLER_22_171 ();
 decap_12 FILLER_22_176 ();
 fill_4 FILLER_22_192 ();
 fill_2 FILLER_22_206 ();
 fill_2 FILLER_22_224 ();
 fill_1 FILLER_22_226 ();
 fill_1 FILLER_22_258 ();
 fill_4 FILLER_22_264 ();
 fill_2 FILLER_22_268 ();
 fill_4 FILLER_22_287 ();
 fill_8 FILLER_22_299 ();
 fill_1 FILLER_22_307 ();
 fill_4 FILLER_22_317 ();
 fill_8 FILLER_22_329 ();
 fill_8 FILLER_22_348 ();
 fill_1 FILLER_22_356 ();
 fill_1 FILLER_22_363 ();
 fill_1 FILLER_22_368 ();
 fill_4 FILLER_22_453 ();
 fill_1 FILLER_22_457 ();
 fill_1 FILLER_22_493 ();
 fill_2 FILLER_22_548 ();
 fill_1 FILLER_22_556 ();
 fill_2 FILLER_22_595 ();
 fill_1 FILLER_22_610 ();
 fill_2 FILLER_22_623 ();
 fill_1 FILLER_22_634 ();
 fill_2 FILLER_22_641 ();
 fill_1 FILLER_22_643 ();
 fill_2 FILLER_22_667 ();
 fill_2 FILLER_22_697 ();
 fill_1 FILLER_22_699 ();
 fill_2 FILLER_22_701 ();
 fill_1 FILLER_22_703 ();
 fill_4 FILLER_22_828 ();
 fill_1 FILLER_22_832 ();
 fill_1 FILLER_22_923 ();
 fill_1 FILLER_22_934 ();
 fill_1 FILLER_22_938 ();
 fill_1 FILLER_22_1008 ();
 fill_1 FILLER_22_1035 ();
 fill_1 FILLER_22_1037 ();
 decap_12 FILLER_23_3 ();
 fill_8 FILLER_23_15 ();
 decap_12 FILLER_23_31 ();
 decap_12 FILLER_23_43 ();
 fill_1 FILLER_23_55 ();
 fill_4 FILLER_23_68 ();
 fill_1 FILLER_23_72 ();
 decap_12 FILLER_23_85 ();
 decap_12 FILLER_23_97 ();
 fill_2 FILLER_23_109 ();
 fill_1 FILLER_23_111 ();
 fill_8 FILLER_23_113 ();
 fill_2 FILLER_23_121 ();
 fill_2 FILLER_23_131 ();
 fill_1 FILLER_23_133 ();
 fill_8 FILLER_23_141 ();
 fill_4 FILLER_23_154 ();
 fill_2 FILLER_23_158 ();
 fill_2 FILLER_23_165 ();
 fill_1 FILLER_23_167 ();
 fill_4 FILLER_23_169 ();
 fill_2 FILLER_23_173 ();
 fill_1 FILLER_23_175 ();
 fill_2 FILLER_23_194 ();
 fill_8 FILLER_23_202 ();
 fill_2 FILLER_23_210 ();
 fill_2 FILLER_23_219 ();
 fill_2 FILLER_23_230 ();
 fill_4 FILLER_23_235 ();
 fill_2 FILLER_23_239 ();
 fill_1 FILLER_23_250 ();
 fill_1 FILLER_23_255 ();
 fill_2 FILLER_23_260 ();
 fill_4 FILLER_23_273 ();
 fill_4 FILLER_23_295 ();
 fill_2 FILLER_23_307 ();
 fill_1 FILLER_23_367 ();
 fill_4 FILLER_23_388 ();
 fill_2 FILLER_23_445 ();
 fill_1 FILLER_23_447 ();
 fill_4 FILLER_23_514 ();
 fill_1 FILLER_23_533 ();
 fill_2 FILLER_23_567 ();
 fill_2 FILLER_23_611 ();
 fill_2 FILLER_23_642 ();
 fill_1 FILLER_23_644 ();
 fill_2 FILLER_23_706 ();
 fill_2 FILLER_23_749 ();
 fill_1 FILLER_23_758 ();
 fill_1 FILLER_23_783 ();
 fill_1 FILLER_23_839 ();
 fill_1 FILLER_23_850 ();
 fill_1 FILLER_23_879 ();
 fill_2 FILLER_23_893 ();
 fill_1 FILLER_23_895 ();
 fill_2 FILLER_23_915 ();
 fill_1 FILLER_23_964 ();
 fill_1 FILLER_23_1007 ();
 fill_1 FILLER_24_3 ();
 fill_4 FILLER_24_22 ();
 fill_2 FILLER_24_26 ();
 fill_1 FILLER_24_34 ();
 fill_4 FILLER_24_50 ();
 fill_1 FILLER_24_61 ();
 fill_2 FILLER_24_72 ();
 fill_1 FILLER_24_83 ();
 fill_2 FILLER_24_85 ();
 fill_4 FILLER_24_99 ();
 fill_4 FILLER_24_110 ();
 fill_2 FILLER_24_114 ();
 fill_1 FILLER_24_116 ();
 fill_8 FILLER_24_125 ();
 fill_2 FILLER_24_133 ();
 fill_1 FILLER_24_135 ();
 fill_1 FILLER_24_157 ();
 decap_12 FILLER_24_173 ();
 fill_8 FILLER_24_185 ();
 fill_2 FILLER_24_193 ();
 fill_1 FILLER_24_195 ();
 fill_4 FILLER_24_207 ();
 fill_2 FILLER_24_221 ();
 fill_1 FILLER_24_229 ();
 fill_8 FILLER_24_242 ();
 fill_2 FILLER_24_250 ();
 fill_4 FILLER_24_260 ();
 fill_1 FILLER_24_264 ();
 fill_1 FILLER_24_268 ();
 fill_2 FILLER_24_290 ();
 fill_1 FILLER_24_292 ();
 fill_1 FILLER_24_298 ();
 fill_1 FILLER_24_307 ();
 fill_4 FILLER_24_309 ();
 fill_2 FILLER_24_313 ();
 fill_1 FILLER_24_315 ();
 fill_2 FILLER_24_319 ();
 fill_1 FILLER_24_321 ();
 fill_4 FILLER_24_329 ();
 fill_2 FILLER_24_333 ();
 fill_2 FILLER_24_365 ();
 fill_2 FILLER_24_408 ();
 fill_1 FILLER_24_419 ();
 fill_4 FILLER_24_446 ();
 fill_1 FILLER_24_450 ();
 fill_2 FILLER_24_471 ();
 fill_1 FILLER_24_477 ();
 fill_1 FILLER_24_494 ();
 fill_1 FILLER_24_504 ();
 fill_2 FILLER_24_517 ();
 fill_4 FILLER_24_528 ();
 fill_1 FILLER_24_553 ();
 fill_1 FILLER_24_587 ();
 fill_1 FILLER_24_607 ();
 fill_1 FILLER_24_658 ();
 fill_4 FILLER_24_696 ();
 fill_2 FILLER_24_715 ();
 fill_2 FILLER_24_737 ();
 fill_1 FILLER_24_747 ();
 fill_1 FILLER_24_755 ();
 fill_2 FILLER_24_813 ();
 fill_2 FILLER_24_846 ();
 fill_2 FILLER_24_869 ();
 fill_4 FILLER_24_918 ();
 fill_2 FILLER_24_922 ();
 fill_1 FILLER_24_951 ();
 fill_2 FILLER_24_957 ();
 fill_1 FILLER_24_981 ();
 fill_1 FILLER_24_1035 ();
 fill_1 FILLER_24_1037 ();
 decap_12 FILLER_25_3 ();
 fill_8 FILLER_25_15 ();
 fill_4 FILLER_25_29 ();
 fill_2 FILLER_25_33 ();
 decap_12 FILLER_25_43 ();
 fill_1 FILLER_25_55 ();
 fill_4 FILLER_25_66 ();
 fill_4 FILLER_25_82 ();
 fill_2 FILLER_25_86 ();
 fill_4 FILLER_25_106 ();
 fill_2 FILLER_25_110 ();
 fill_1 FILLER_25_133 ();
 fill_8 FILLER_25_143 ();
 fill_4 FILLER_25_159 ();
 fill_1 FILLER_25_163 ();
 fill_1 FILLER_25_167 ();
 fill_4 FILLER_25_169 ();
 fill_1 FILLER_25_173 ();
 fill_4 FILLER_25_179 ();
 fill_1 FILLER_25_223 ();
 fill_2 FILLER_25_233 ();
 fill_1 FILLER_25_281 ();
 fill_1 FILLER_25_310 ();
 fill_2 FILLER_25_318 ();
 decap_12 FILLER_25_346 ();
 fill_1 FILLER_25_358 ();
 fill_1 FILLER_25_372 ();
 fill_1 FILLER_25_376 ();
 fill_2 FILLER_25_390 ();
 fill_1 FILLER_25_406 ();
 fill_1 FILLER_25_412 ();
 fill_2 FILLER_25_446 ();
 fill_2 FILLER_25_461 ();
 fill_1 FILLER_25_483 ();
 fill_2 FILLER_25_512 ();
 fill_4 FILLER_25_534 ();
 fill_1 FILLER_25_559 ();
 fill_1 FILLER_25_579 ();
 fill_1 FILLER_25_606 ();
 fill_1 FILLER_25_626 ();
 fill_1 FILLER_25_636 ();
 fill_1 FILLER_25_646 ();
 fill_4 FILLER_25_660 ();
 fill_1 FILLER_25_664 ();
 fill_4 FILLER_25_704 ();
 fill_1 FILLER_25_721 ();
 fill_1 FILLER_25_749 ();
 fill_1 FILLER_25_763 ();
 fill_1 FILLER_25_783 ();
 fill_1 FILLER_25_821 ();
 fill_1 FILLER_25_846 ();
 fill_4 FILLER_25_897 ();
 fill_1 FILLER_25_901 ();
 fill_2 FILLER_25_908 ();
 fill_1 FILLER_25_910 ();
 fill_1 FILLER_25_940 ();
 fill_2 FILLER_25_950 ();
 fill_1 FILLER_25_1037 ();
 fill_4 FILLER_26_3 ();
 fill_2 FILLER_26_7 ();
 fill_4 FILLER_26_23 ();
 fill_1 FILLER_26_27 ();
 fill_4 FILLER_26_50 ();
 fill_2 FILLER_26_54 ();
 fill_4 FILLER_26_59 ();
 fill_2 FILLER_26_63 ();
 fill_8 FILLER_26_100 ();
 fill_1 FILLER_26_108 ();
 fill_4 FILLER_26_114 ();
 fill_1 FILLER_26_118 ();
 fill_2 FILLER_26_129 ();
 fill_1 FILLER_26_131 ();
 fill_2 FILLER_26_148 ();
 fill_1 FILLER_26_150 ();
 fill_4 FILLER_26_154 ();
 fill_2 FILLER_26_158 ();
 fill_1 FILLER_26_160 ();
 fill_1 FILLER_26_179 ();
 fill_1 FILLER_26_214 ();
 fill_4 FILLER_26_238 ();
 fill_1 FILLER_26_242 ();
 fill_4 FILLER_26_248 ();
 fill_4 FILLER_26_253 ();
 fill_8 FILLER_26_262 ();
 fill_4 FILLER_26_295 ();
 fill_2 FILLER_26_299 ();
 fill_1 FILLER_26_301 ();
 fill_2 FILLER_26_309 ();
 fill_2 FILLER_26_332 ();
 fill_2 FILLER_26_398 ();
 fill_2 FILLER_26_412 ();
 fill_2 FILLER_26_418 ();
 fill_2 FILLER_26_442 ();
 fill_4 FILLER_26_503 ();
 fill_1 FILLER_26_514 ();
 decap_12 FILLER_26_518 ();
 fill_2 FILLER_26_530 ();
 fill_2 FILLER_26_562 ();
 fill_2 FILLER_26_592 ();
 fill_1 FILLER_26_643 ();
 fill_4 FILLER_26_668 ();
 fill_4 FILLER_26_676 ();
 fill_1 FILLER_26_680 ();
 fill_2 FILLER_26_701 ();
 fill_2 FILLER_26_730 ();
 fill_2 FILLER_26_745 ();
 fill_1 FILLER_26_747 ();
 fill_1 FILLER_26_755 ();
 fill_2 FILLER_26_757 ();
 fill_1 FILLER_26_759 ();
 fill_4 FILLER_26_780 ();
 fill_1 FILLER_26_784 ();
 fill_2 FILLER_26_794 ();
 fill_1 FILLER_26_811 ();
 fill_1 FILLER_26_848 ();
 fill_1 FILLER_26_858 ();
 fill_1 FILLER_26_872 ();
 fill_2 FILLER_26_902 ();
 fill_1 FILLER_26_923 ();
 fill_8 FILLER_26_934 ();
 fill_1 FILLER_26_942 ();
 fill_2 FILLER_26_964 ();
 fill_2 FILLER_26_975 ();
 fill_1 FILLER_26_987 ();
 fill_1 FILLER_26_1009 ();
 fill_1 FILLER_26_1031 ();
 fill_1 FILLER_26_1035 ();
 fill_1 FILLER_26_1037 ();
 decap_12 FILLER_27_3 ();
 decap_12 FILLER_27_15 ();
 fill_4 FILLER_27_27 ();
 fill_4 FILLER_27_39 ();
 fill_2 FILLER_27_54 ();
 fill_1 FILLER_27_62 ();
 fill_4 FILLER_27_66 ();
 fill_1 FILLER_27_87 ();
 fill_8 FILLER_27_91 ();
 fill_1 FILLER_27_99 ();
 decap_12 FILLER_27_127 ();
 fill_8 FILLER_27_139 ();
 fill_1 FILLER_27_147 ();
 fill_8 FILLER_27_160 ();
 fill_4 FILLER_27_169 ();
 fill_1 FILLER_27_173 ();
 fill_1 FILLER_27_186 ();
 fill_1 FILLER_27_197 ();
 fill_1 FILLER_27_245 ();
 fill_1 FILLER_27_267 ();
 fill_4 FILLER_27_276 ();
 fill_4 FILLER_27_314 ();
 fill_2 FILLER_27_318 ();
 fill_4 FILLER_27_324 ();
 fill_2 FILLER_27_328 ();
 fill_1 FILLER_27_330 ();
 fill_2 FILLER_27_334 ();
 fill_2 FILLER_27_337 ();
 fill_1 FILLER_27_348 ();
 fill_1 FILLER_27_375 ();
 fill_2 FILLER_27_390 ();
 fill_4 FILLER_27_393 ();
 fill_2 FILLER_27_397 ();
 fill_1 FILLER_27_407 ();
 fill_2 FILLER_27_416 ();
 fill_2 FILLER_27_439 ();
 fill_1 FILLER_27_441 ();
 fill_2 FILLER_27_469 ();
 fill_1 FILLER_27_503 ();
 fill_1 FILLER_27_505 ();
 fill_8 FILLER_27_529 ();
 fill_2 FILLER_27_537 ();
 fill_2 FILLER_27_545 ();
 fill_8 FILLER_27_550 ();
 fill_2 FILLER_27_558 ();
 fill_1 FILLER_27_561 ();
 fill_4 FILLER_27_571 ();
 fill_2 FILLER_27_613 ();
 fill_1 FILLER_27_615 ();
 fill_8 FILLER_27_617 ();
 fill_1 FILLER_27_625 ();
 fill_1 FILLER_27_652 ();
 fill_1 FILLER_27_671 ();
 fill_2 FILLER_27_679 ();
 fill_1 FILLER_27_707 ();
 fill_1 FILLER_27_737 ();
 fill_4 FILLER_27_760 ();
 fill_1 FILLER_27_764 ();
 fill_1 FILLER_27_783 ();
 fill_1 FILLER_27_876 ();
 fill_1 FILLER_27_887 ();
 fill_1 FILLER_27_895 ();
 fill_2 FILLER_27_906 ();
 fill_4 FILLER_27_931 ();
 fill_2 FILLER_27_935 ();
 fill_1 FILLER_27_937 ();
 fill_2 FILLER_27_944 ();
 fill_2 FILLER_27_962 ();
 fill_1 FILLER_27_1002 ();
 fill_2 FILLER_27_1015 ();
 fill_1 FILLER_27_1037 ();
 fill_2 FILLER_28_3 ();
 fill_4 FILLER_28_12 ();
 fill_2 FILLER_28_16 ();
 fill_4 FILLER_28_24 ();
 fill_2 FILLER_28_34 ();
 fill_8 FILLER_28_40 ();
 fill_2 FILLER_28_48 ();
 fill_1 FILLER_28_50 ();
 fill_2 FILLER_28_69 ();
 fill_1 FILLER_28_71 ();
 fill_8 FILLER_28_75 ();
 fill_1 FILLER_28_83 ();
 fill_4 FILLER_28_107 ();
 fill_4 FILLER_28_136 ();
 fill_4 FILLER_28_146 ();
 fill_1 FILLER_28_150 ();
 decap_12 FILLER_28_157 ();
 fill_1 FILLER_28_197 ();
 fill_2 FILLER_28_211 ();
 fill_1 FILLER_28_251 ();
 fill_4 FILLER_28_264 ();
 fill_1 FILLER_28_268 ();
 fill_4 FILLER_28_277 ();
 fill_2 FILLER_28_281 ();
 fill_8 FILLER_28_289 ();
 fill_4 FILLER_28_301 ();
 fill_2 FILLER_28_305 ();
 fill_1 FILLER_28_307 ();
 fill_4 FILLER_28_309 ();
 fill_1 FILLER_28_313 ();
 fill_4 FILLER_28_339 ();
 fill_1 FILLER_28_343 ();
 fill_8 FILLER_28_371 ();
 fill_2 FILLER_28_399 ();
 fill_1 FILLER_28_401 ();
 fill_1 FILLER_28_405 ();
 fill_2 FILLER_28_418 ();
 fill_2 FILLER_28_441 ();
 fill_2 FILLER_28_449 ();
 fill_1 FILLER_28_477 ();
 fill_1 FILLER_28_488 ();
 fill_4 FILLER_28_501 ();
 fill_2 FILLER_28_510 ();
 fill_1 FILLER_28_540 ();
 fill_2 FILLER_28_550 ();
 fill_1 FILLER_28_552 ();
 fill_4 FILLER_28_573 ();
 fill_1 FILLER_28_577 ();
 fill_1 FILLER_28_584 ();
 fill_2 FILLER_28_618 ();
 fill_2 FILLER_28_641 ();
 fill_1 FILLER_28_643 ();
 fill_1 FILLER_28_699 ();
 fill_1 FILLER_28_737 ();
 fill_2 FILLER_28_747 ();
 fill_1 FILLER_28_780 ();
 fill_1 FILLER_28_799 ();
 fill_1 FILLER_28_806 ();
 fill_1 FILLER_28_813 ();
 fill_4 FILLER_28_881 ();
 fill_2 FILLER_28_885 ();
 fill_4 FILLER_28_902 ();
 fill_4 FILLER_28_920 ();
 fill_2 FILLER_28_954 ();
 fill_1 FILLER_28_976 ();
 fill_2 FILLER_28_1031 ();
 fill_1 FILLER_28_1037 ();
 fill_4 FILLER_29_3 ();
 fill_1 FILLER_29_7 ();
 decap_12 FILLER_29_13 ();
 fill_2 FILLER_29_25 ();
 fill_2 FILLER_29_31 ();
 fill_4 FILLER_29_51 ();
 fill_1 FILLER_29_55 ();
 fill_1 FILLER_29_65 ();
 fill_1 FILLER_29_72 ();
 fill_2 FILLER_29_86 ();
 fill_2 FILLER_29_109 ();
 fill_1 FILLER_29_111 ();
 decap_12 FILLER_29_126 ();
 fill_1 FILLER_29_138 ();
 fill_4 FILLER_29_147 ();
 fill_2 FILLER_29_206 ();
 fill_1 FILLER_29_223 ();
 fill_1 FILLER_29_264 ();
 fill_2 FILLER_29_274 ();
 fill_2 FILLER_29_297 ();
 fill_1 FILLER_29_299 ();
 fill_2 FILLER_29_320 ();
 fill_4 FILLER_29_332 ();
 fill_2 FILLER_29_344 ();
 fill_1 FILLER_29_346 ();
 fill_2 FILLER_29_367 ();
 fill_1 FILLER_29_377 ();
 fill_4 FILLER_29_384 ();
 fill_2 FILLER_29_431 ();
 fill_1 FILLER_29_433 ();
 fill_4 FILLER_29_460 ();
 fill_1 FILLER_29_464 ();
 fill_1 FILLER_29_498 ();
 fill_2 FILLER_29_531 ();
 fill_1 FILLER_29_533 ();
 fill_2 FILLER_29_609 ();
 fill_1 FILLER_29_625 ();
 fill_2 FILLER_29_670 ();
 fill_1 FILLER_29_682 ();
 fill_2 FILLER_29_697 ();
 fill_1 FILLER_29_727 ();
 fill_2 FILLER_29_729 ();
 fill_1 FILLER_29_783 ();
 fill_1 FILLER_29_833 ();
 fill_2 FILLER_29_841 ();
 fill_1 FILLER_29_843 ();
 fill_2 FILLER_29_864 ();
 fill_1 FILLER_29_875 ();
 fill_2 FILLER_29_897 ();
 fill_1 FILLER_29_899 ();
 fill_2 FILLER_29_923 ();
 fill_1 FILLER_29_925 ();
 fill_2 FILLER_29_935 ();
 fill_1 FILLER_29_962 ();
 fill_2 FILLER_30_3 ();
 fill_1 FILLER_30_5 ();
 fill_8 FILLER_30_12 ();
 decap_12 FILLER_30_38 ();
 decap_12 FILLER_30_50 ();
 fill_4 FILLER_30_62 ();
 fill_2 FILLER_30_66 ();
 fill_1 FILLER_30_68 ();
 fill_2 FILLER_30_88 ();
 fill_4 FILLER_30_109 ();
 fill_1 FILLER_30_113 ();
 fill_8 FILLER_30_118 ();
 fill_1 FILLER_30_139 ();
 decap_12 FILLER_30_145 ();
 fill_8 FILLER_30_157 ();
 fill_2 FILLER_30_170 ();
 fill_1 FILLER_30_172 ();
 fill_1 FILLER_30_195 ();
 fill_2 FILLER_30_249 ();
 fill_1 FILLER_30_251 ();
 fill_8 FILLER_30_257 ();
 fill_2 FILLER_30_265 ();
 fill_2 FILLER_30_278 ();
 fill_1 FILLER_30_280 ();
 fill_2 FILLER_30_292 ();
 fill_8 FILLER_30_297 ();
 fill_2 FILLER_30_305 ();
 fill_1 FILLER_30_307 ();
 fill_4 FILLER_30_309 ();
 fill_1 FILLER_30_313 ();
 fill_2 FILLER_30_319 ();
 fill_1 FILLER_30_321 ();
 fill_8 FILLER_30_356 ();
 fill_1 FILLER_30_370 ();
 fill_4 FILLER_30_391 ();
 fill_4 FILLER_30_415 ();
 fill_1 FILLER_30_419 ();
 fill_8 FILLER_30_421 ();
 fill_2 FILLER_30_429 ();
 fill_1 FILLER_30_431 ();
 fill_1 FILLER_30_475 ();
 fill_2 FILLER_30_498 ();
 fill_1 FILLER_30_500 ();
 fill_1 FILLER_30_511 ();
 fill_4 FILLER_30_539 ();
 fill_2 FILLER_30_552 ();
 fill_4 FILLER_30_581 ();
 fill_2 FILLER_30_585 ();
 fill_1 FILLER_30_587 ();
 fill_4 FILLER_30_598 ();
 fill_1 FILLER_30_602 ();
 fill_2 FILLER_30_613 ();
 fill_1 FILLER_30_631 ();
 fill_2 FILLER_30_641 ();
 fill_1 FILLER_30_643 ();
 fill_2 FILLER_30_645 ();
 fill_1 FILLER_30_659 ();
 fill_4 FILLER_30_680 ();
 fill_1 FILLER_30_699 ();
 fill_1 FILLER_30_701 ();
 fill_1 FILLER_30_717 ();
 fill_1 FILLER_30_764 ();
 fill_2 FILLER_30_787 ();
 fill_1 FILLER_30_834 ();
 fill_1 FILLER_30_843 ();
 fill_2 FILLER_30_878 ();
 fill_1 FILLER_30_880 ();
 fill_2 FILLER_30_890 ();
 fill_1 FILLER_30_892 ();
 fill_1 FILLER_30_917 ();
 fill_2 FILLER_30_965 ();
 fill_1 FILLER_30_979 ();
 fill_2 FILLER_30_1025 ();
 fill_1 FILLER_30_1037 ();
 fill_4 FILLER_31_3 ();
 decap_12 FILLER_31_17 ();
 fill_1 FILLER_31_29 ();
 fill_8 FILLER_31_37 ();
 fill_2 FILLER_31_45 ();
 fill_2 FILLER_31_54 ();
 fill_2 FILLER_31_64 ();
 fill_1 FILLER_31_66 ();
 fill_2 FILLER_31_74 ();
 fill_1 FILLER_31_81 ();
 fill_2 FILLER_31_110 ();
 fill_4 FILLER_31_119 ();
 fill_2 FILLER_31_152 ();
 fill_1 FILLER_31_154 ();
 fill_4 FILLER_31_192 ();
 fill_2 FILLER_31_209 ();
 fill_1 FILLER_31_211 ();
 fill_2 FILLER_31_271 ();
 fill_2 FILLER_31_285 ();
 fill_1 FILLER_31_287 ();
 fill_2 FILLER_31_325 ();
 fill_2 FILLER_31_334 ();
 fill_4 FILLER_31_337 ();
 fill_1 FILLER_31_341 ();
 fill_4 FILLER_31_349 ();
 decap_12 FILLER_31_374 ();
 fill_4 FILLER_31_386 ();
 fill_2 FILLER_31_390 ();
 fill_4 FILLER_31_416 ();
 fill_1 FILLER_31_447 ();
 fill_4 FILLER_31_449 ();
 fill_2 FILLER_31_453 ();
 fill_2 FILLER_31_460 ();
 fill_1 FILLER_31_503 ();
 fill_1 FILLER_31_534 ();
 fill_2 FILLER_31_558 ();
 fill_8 FILLER_31_561 ();
 fill_1 FILLER_31_569 ();
 fill_4 FILLER_31_579 ();
 fill_1 FILLER_31_598 ();
 fill_4 FILLER_31_665 ();
 fill_1 FILLER_31_673 ();
 fill_1 FILLER_31_727 ();
 fill_1 FILLER_31_748 ();
 fill_1 FILLER_31_759 ();
 fill_1 FILLER_31_780 ();
 fill_1 FILLER_31_797 ();
 fill_1 FILLER_31_830 ();
 fill_1 FILLER_31_847 ();
 fill_1 FILLER_31_857 ();
 fill_2 FILLER_31_870 ();
 fill_4 FILLER_31_892 ();
 fill_2 FILLER_31_935 ();
 fill_4 FILLER_31_940 ();
 fill_4 FILLER_31_980 ();
 fill_1 FILLER_31_984 ();
 fill_1 FILLER_31_994 ();
 fill_1 FILLER_32_3 ();
 fill_4 FILLER_32_24 ();
 fill_1 FILLER_32_29 ();
 fill_2 FILLER_32_37 ();
 fill_1 FILLER_32_39 ();
 fill_2 FILLER_32_54 ();
 fill_1 FILLER_32_56 ();
 fill_8 FILLER_32_103 ();
 fill_1 FILLER_32_111 ();
 fill_4 FILLER_32_136 ();
 fill_2 FILLER_32_141 ();
 fill_2 FILLER_32_207 ();
 fill_1 FILLER_32_209 ();
 fill_1 FILLER_32_232 ();
 fill_1 FILLER_32_251 ();
 fill_2 FILLER_32_253 ();
 fill_1 FILLER_32_270 ();
 fill_4 FILLER_32_287 ();
 fill_1 FILLER_32_291 ();
 fill_4 FILLER_32_303 ();
 fill_1 FILLER_32_307 ();
 fill_1 FILLER_32_309 ();
 fill_1 FILLER_32_320 ();
 fill_1 FILLER_32_337 ();
 fill_2 FILLER_32_362 ();
 fill_2 FILLER_32_392 ();
 fill_1 FILLER_32_394 ();
 fill_1 FILLER_32_421 ();
 fill_2 FILLER_32_433 ();
 fill_1 FILLER_32_449 ();
 fill_4 FILLER_32_470 ();
 fill_2 FILLER_32_474 ();
 fill_8 FILLER_32_483 ();
 fill_1 FILLER_32_517 ();
 fill_1 FILLER_32_526 ();
 fill_4 FILLER_32_551 ();
 fill_1 FILLER_32_555 ();
 fill_2 FILLER_32_585 ();
 fill_1 FILLER_32_587 ();
 fill_2 FILLER_32_610 ();
 fill_1 FILLER_32_612 ();
 fill_1 FILLER_32_639 ();
 fill_4 FILLER_32_657 ();
 fill_1 FILLER_32_661 ();
 fill_1 FILLER_32_686 ();
 fill_1 FILLER_32_727 ();
 fill_1 FILLER_32_741 ();
 fill_1 FILLER_32_751 ();
 fill_1 FILLER_32_771 ();
 fill_2 FILLER_32_813 ();
 fill_4 FILLER_32_863 ();
 fill_1 FILLER_32_867 ();
 fill_4 FILLER_32_869 ();
 fill_2 FILLER_32_873 ();
 fill_1 FILLER_32_875 ();
 fill_1 FILLER_32_896 ();
 fill_1 FILLER_32_934 ();
 fill_1 FILLER_32_962 ();
 fill_2 FILLER_32_978 ();
 fill_1 FILLER_32_993 ();
 fill_1 FILLER_32_1037 ();
 fill_2 FILLER_33_23 ();
 fill_4 FILLER_33_36 ();
 fill_2 FILLER_33_40 ();
 fill_8 FILLER_33_45 ();
 fill_2 FILLER_33_53 ();
 fill_1 FILLER_33_55 ();
 fill_2 FILLER_33_57 ();
 fill_1 FILLER_33_59 ();
 fill_4 FILLER_33_63 ();
 fill_2 FILLER_33_67 ();
 fill_1 FILLER_33_78 ();
 fill_2 FILLER_33_113 ();
 fill_1 FILLER_33_115 ();
 fill_4 FILLER_33_136 ();
 fill_4 FILLER_33_150 ();
 fill_2 FILLER_33_154 ();
 fill_1 FILLER_33_156 ();
 fill_2 FILLER_33_178 ();
 fill_1 FILLER_33_180 ();
 fill_2 FILLER_33_193 ();
 fill_1 FILLER_33_195 ();
 fill_2 FILLER_33_221 ();
 fill_1 FILLER_33_223 ();
 fill_1 FILLER_33_242 ();
 fill_8 FILLER_33_246 ();
 fill_2 FILLER_33_254 ();
 fill_8 FILLER_33_263 ();
 fill_2 FILLER_33_278 ();
 fill_1 FILLER_33_284 ();
 fill_2 FILLER_33_299 ();
 fill_2 FILLER_33_305 ();
 fill_1 FILLER_33_307 ();
 fill_2 FILLER_33_315 ();
 fill_4 FILLER_33_332 ();
 fill_4 FILLER_33_352 ();
 fill_2 FILLER_33_356 ();
 fill_1 FILLER_33_374 ();
 fill_2 FILLER_33_401 ();
 fill_4 FILLER_33_473 ();
 fill_2 FILLER_33_477 ();
 fill_1 FILLER_33_479 ();
 fill_2 FILLER_33_502 ();
 fill_2 FILLER_33_505 ();
 fill_1 FILLER_33_507 ();
 fill_2 FILLER_33_523 ();
 fill_1 FILLER_33_525 ();
 decap_12 FILLER_33_566 ();
 fill_8 FILLER_33_587 ();
 fill_1 FILLER_33_595 ();
 fill_1 FILLER_33_605 ();
 fill_4 FILLER_33_612 ();
 fill_4 FILLER_33_624 ();
 fill_4 FILLER_33_637 ();
 fill_1 FILLER_33_641 ();
 fill_2 FILLER_33_654 ();
 fill_1 FILLER_33_659 ();
 fill_1 FILLER_33_749 ();
 fill_2 FILLER_33_800 ();
 fill_1 FILLER_33_839 ();
 fill_4 FILLER_33_844 ();
 fill_1 FILLER_33_848 ();
 fill_1 FILLER_33_858 ();
 fill_2 FILLER_33_953 ();
 fill_2 FILLER_33_978 ();
 fill_2 FILLER_33_1006 ();
 fill_2 FILLER_33_1009 ();
 fill_4 FILLER_34_3 ();
 fill_1 FILLER_34_7 ();
 fill_2 FILLER_34_52 ();
 fill_2 FILLER_34_82 ();
 fill_1 FILLER_34_128 ();
 fill_2 FILLER_34_138 ();
 fill_1 FILLER_34_185 ();
 fill_2 FILLER_34_194 ();
 fill_2 FILLER_34_222 ();
 fill_2 FILLER_34_231 ();
 fill_1 FILLER_34_233 ();
 fill_2 FILLER_34_245 ();
 fill_1 FILLER_34_247 ();
 fill_4 FILLER_34_260 ();
 fill_2 FILLER_34_264 ();
 fill_1 FILLER_34_266 ();
 fill_2 FILLER_34_306 ();
 fill_1 FILLER_34_331 ();
 fill_1 FILLER_34_346 ();
 fill_2 FILLER_34_355 ();
 fill_1 FILLER_34_369 ();
 fill_8 FILLER_34_410 ();
 fill_2 FILLER_34_418 ();
 fill_1 FILLER_34_421 ();
 fill_4 FILLER_34_435 ();
 fill_4 FILLER_34_444 ();
 fill_2 FILLER_34_466 ();
 fill_1 FILLER_34_468 ();
 fill_8 FILLER_34_500 ();
 fill_1 FILLER_34_508 ();
 fill_2 FILLER_34_530 ();
 fill_2 FILLER_34_533 ();
 fill_1 FILLER_34_535 ();
 fill_2 FILLER_34_557 ();
 fill_1 FILLER_34_559 ();
 fill_1 FILLER_34_595 ();
 fill_2 FILLER_34_642 ();
 fill_1 FILLER_34_679 ();
 fill_1 FILLER_34_725 ();
 fill_2 FILLER_34_757 ();
 fill_1 FILLER_34_788 ();
 fill_2 FILLER_34_810 ();
 fill_1 FILLER_34_864 ();
 fill_2 FILLER_34_921 ();
 fill_1 FILLER_34_923 ();
 fill_8 FILLER_34_925 ();
 fill_1 FILLER_34_933 ();
 fill_1 FILLER_34_979 ();
 fill_1 FILLER_34_1037 ();
 decap_12 FILLER_35_6 ();
 fill_2 FILLER_35_18 ();
 fill_2 FILLER_35_71 ();
 fill_4 FILLER_35_76 ();
 fill_2 FILLER_35_80 ();
 fill_2 FILLER_35_110 ();
 fill_2 FILLER_35_155 ();
 fill_1 FILLER_35_157 ();
 fill_2 FILLER_35_169 ();
 fill_2 FILLER_35_176 ();
 fill_1 FILLER_35_223 ();
 fill_2 FILLER_35_225 ();
 fill_1 FILLER_35_227 ();
 fill_1 FILLER_35_241 ();
 fill_1 FILLER_35_255 ();
 fill_4 FILLER_35_281 ();
 fill_1 FILLER_35_285 ();
 fill_1 FILLER_35_307 ();
 fill_2 FILLER_35_316 ();
 fill_4 FILLER_35_331 ();
 fill_1 FILLER_35_335 ();
 fill_2 FILLER_35_352 ();
 fill_1 FILLER_35_373 ();
 fill_2 FILLER_35_382 ();
 fill_1 FILLER_35_384 ();
 fill_1 FILLER_35_403 ();
 fill_2 FILLER_35_446 ();
 fill_2 FILLER_35_456 ();
 fill_4 FILLER_35_483 ();
 fill_1 FILLER_35_487 ();
 fill_4 FILLER_35_505 ();
 fill_1 FILLER_35_509 ();
 decap_12 FILLER_35_548 ();
 fill_1 FILLER_35_582 ();
 fill_4 FILLER_35_591 ();
 fill_2 FILLER_35_599 ();
 fill_1 FILLER_35_601 ();
 fill_4 FILLER_35_609 ();
 fill_2 FILLER_35_613 ();
 fill_1 FILLER_35_615 ();
 fill_4 FILLER_35_637 ();
 fill_2 FILLER_35_641 ();
 fill_1 FILLER_35_643 ();
 fill_2 FILLER_35_650 ();
 fill_1 FILLER_35_733 ();
 fill_1 FILLER_35_754 ();
 fill_2 FILLER_35_782 ();
 fill_2 FILLER_35_824 ();
 fill_1 FILLER_35_826 ();
 fill_1 FILLER_35_839 ();
 fill_8 FILLER_35_841 ();
 fill_1 FILLER_35_849 ();
 fill_1 FILLER_35_885 ();
 fill_1 FILLER_35_895 ();
 fill_1 FILLER_35_897 ();
 fill_2 FILLER_35_913 ();
 fill_4 FILLER_35_944 ();
 fill_1 FILLER_35_948 ();
 fill_1 FILLER_35_966 ();
 fill_2 FILLER_35_1005 ();
 fill_1 FILLER_35_1007 ();
 decap_12 FILLER_36_3 ();
 decap_12 FILLER_36_15 ();
 fill_1 FILLER_36_27 ();
 fill_1 FILLER_36_67 ();
 fill_4 FILLER_36_77 ();
 fill_2 FILLER_36_81 ();
 fill_1 FILLER_36_83 ();
 fill_1 FILLER_36_105 ();
 fill_1 FILLER_36_125 ();
 fill_4 FILLER_36_135 ();
 fill_1 FILLER_36_139 ();
 fill_4 FILLER_36_141 ();
 fill_2 FILLER_36_145 ();
 fill_4 FILLER_36_166 ();
 fill_2 FILLER_36_200 ();
 fill_1 FILLER_36_202 ();
 fill_1 FILLER_36_218 ();
 fill_2 FILLER_36_250 ();
 fill_4 FILLER_36_253 ();
 fill_1 FILLER_36_277 ();
 fill_4 FILLER_36_283 ();
 fill_2 FILLER_36_287 ();
 fill_4 FILLER_36_302 ();
 fill_2 FILLER_36_306 ();
 fill_1 FILLER_36_324 ();
 fill_2 FILLER_36_329 ();
 fill_1 FILLER_36_331 ();
 fill_1 FILLER_36_349 ();
 fill_2 FILLER_36_354 ();
 fill_8 FILLER_36_365 ();
 fill_2 FILLER_36_387 ();
 fill_1 FILLER_36_389 ();
 fill_4 FILLER_36_415 ();
 fill_1 FILLER_36_419 ();
 fill_2 FILLER_36_421 ();
 fill_1 FILLER_36_423 ();
 fill_1 FILLER_36_430 ();
 fill_1 FILLER_36_446 ();
 fill_1 FILLER_36_475 ();
 fill_1 FILLER_36_477 ();
 fill_4 FILLER_36_526 ();
 fill_2 FILLER_36_530 ();
 fill_4 FILLER_36_533 ();
 fill_1 FILLER_36_537 ();
 fill_4 FILLER_36_582 ();
 fill_2 FILLER_36_586 ();
 fill_2 FILLER_36_589 ();
 fill_1 FILLER_36_591 ();
 fill_8 FILLER_36_613 ();
 fill_1 FILLER_36_710 ();
 fill_2 FILLER_36_741 ();
 fill_1 FILLER_36_795 ();
 fill_1 FILLER_36_811 ();
 fill_2 FILLER_36_839 ();
 fill_2 FILLER_36_860 ();
 fill_2 FILLER_36_921 ();
 fill_1 FILLER_36_923 ();
 fill_1 FILLER_36_934 ();
 fill_2 FILLER_36_947 ();
 fill_1 FILLER_36_999 ();
 fill_1 FILLER_36_1015 ();
 fill_1 FILLER_36_1037 ();
 decap_12 FILLER_37_3 ();
 fill_2 FILLER_37_15 ();
 fill_8 FILLER_37_46 ();
 fill_2 FILLER_37_54 ();
 fill_1 FILLER_37_100 ();
 fill_1 FILLER_37_116 ();
 fill_8 FILLER_37_134 ();
 fill_1 FILLER_37_142 ();
 fill_1 FILLER_37_151 ();
 fill_8 FILLER_37_193 ();
 fill_1 FILLER_37_201 ();
 fill_2 FILLER_37_221 ();
 fill_1 FILLER_37_223 ();
 fill_2 FILLER_37_232 ();
 fill_2 FILLER_37_288 ();
 fill_2 FILLER_37_334 ();
 fill_4 FILLER_37_337 ();
 fill_2 FILLER_37_341 ();
 fill_1 FILLER_37_343 ();
 fill_2 FILLER_37_351 ();
 fill_1 FILLER_37_353 ();
 fill_2 FILLER_37_372 ();
 fill_1 FILLER_37_374 ();
 fill_8 FILLER_37_383 ();
 fill_1 FILLER_37_391 ();
 fill_2 FILLER_37_393 ();
 fill_2 FILLER_37_446 ();
 decap_12 FILLER_37_478 ();
 decap_12 FILLER_37_490 ();
 fill_2 FILLER_37_502 ();
 fill_2 FILLER_37_525 ();
 fill_1 FILLER_37_527 ();
 fill_4 FILLER_37_554 ();
 fill_2 FILLER_37_558 ();
 fill_2 FILLER_37_564 ();
 fill_4 FILLER_37_617 ();
 fill_1 FILLER_37_621 ();
 fill_4 FILLER_37_630 ();
 fill_2 FILLER_37_664 ();
 fill_1 FILLER_37_666 ();
 fill_1 FILLER_37_720 ();
 fill_1 FILLER_37_727 ();
 fill_2 FILLER_37_768 ();
 fill_1 FILLER_37_783 ();
 fill_1 FILLER_37_789 ();
 fill_1 FILLER_37_799 ();
 fill_1 FILLER_37_867 ();
 fill_1 FILLER_37_895 ();
 fill_1 FILLER_37_919 ();
 fill_1 FILLER_37_987 ();
 fill_1 FILLER_37_1018 ();
 fill_4 FILLER_37_1034 ();
 decap_12 FILLER_38_3 ();
 fill_8 FILLER_38_15 ();
 fill_1 FILLER_38_23 ();
 fill_1 FILLER_38_27 ();
 fill_4 FILLER_38_64 ();
 fill_8 FILLER_38_85 ();
 fill_1 FILLER_38_93 ();
 fill_1 FILLER_38_119 ();
 fill_1 FILLER_38_127 ();
 fill_8 FILLER_38_162 ();
 fill_2 FILLER_38_170 ();
 fill_1 FILLER_38_172 ();
 fill_2 FILLER_38_249 ();
 fill_1 FILLER_38_251 ();
 fill_4 FILLER_38_262 ();
 fill_2 FILLER_38_266 ();
 fill_2 FILLER_38_276 ();
 fill_4 FILLER_38_281 ();
 fill_2 FILLER_38_285 ();
 fill_1 FILLER_38_287 ();
 fill_1 FILLER_38_297 ();
 fill_1 FILLER_38_307 ();
 fill_4 FILLER_38_315 ();
 fill_2 FILLER_38_319 ();
 fill_1 FILLER_38_321 ();
 fill_8 FILLER_38_326 ();
 fill_2 FILLER_38_334 ();
 fill_1 FILLER_38_336 ();
 decap_12 FILLER_38_352 ();
 fill_4 FILLER_38_373 ();
 fill_2 FILLER_38_377 ();
 fill_8 FILLER_38_390 ();
 fill_2 FILLER_38_398 ();
 fill_1 FILLER_38_400 ();
 fill_2 FILLER_38_418 ();
 fill_1 FILLER_38_421 ();
 fill_1 FILLER_38_428 ();
 fill_2 FILLER_38_443 ();
 fill_1 FILLER_38_450 ();
 fill_4 FILLER_38_471 ();
 fill_1 FILLER_38_475 ();
 decap_12 FILLER_38_520 ();
 fill_2 FILLER_38_537 ();
 fill_4 FILLER_38_547 ();
 fill_2 FILLER_38_578 ();
 fill_1 FILLER_38_580 ();
 fill_2 FILLER_38_663 ();
 fill_1 FILLER_38_693 ();
 fill_1 FILLER_38_744 ();
 fill_2 FILLER_38_754 ();
 fill_1 FILLER_38_761 ();
 fill_1 FILLER_38_771 ();
 fill_1 FILLER_38_811 ();
 fill_1 FILLER_38_867 ();
 fill_1 FILLER_38_869 ();
 fill_2 FILLER_38_880 ();
 fill_1 FILLER_38_891 ();
 fill_2 FILLER_38_912 ();
 fill_2 FILLER_38_981 ();
 fill_2 FILLER_38_1012 ();
 fill_2 FILLER_38_1034 ();
 fill_1 FILLER_38_1037 ();
 decap_12 FILLER_39_3 ();
 decap_12 FILLER_39_15 ();
 fill_4 FILLER_39_27 ();
 fill_1 FILLER_39_31 ();
 fill_2 FILLER_39_40 ();
 fill_1 FILLER_39_42 ();
 fill_1 FILLER_39_55 ();
 fill_4 FILLER_39_57 ();
 fill_1 FILLER_39_61 ();
 fill_2 FILLER_39_104 ();
 fill_1 FILLER_39_106 ();
 fill_4 FILLER_39_113 ();
 fill_2 FILLER_39_117 ();
 fill_1 FILLER_39_119 ();
 fill_2 FILLER_39_136 ();
 fill_1 FILLER_39_138 ();
 fill_4 FILLER_39_149 ();
 fill_1 FILLER_39_163 ();
 fill_2 FILLER_39_169 ();
 fill_1 FILLER_39_171 ();
 fill_2 FILLER_39_206 ();
 fill_1 FILLER_39_208 ();
 fill_1 FILLER_39_213 ();
 fill_4 FILLER_39_238 ();
 fill_1 FILLER_39_247 ();
 fill_2 FILLER_39_273 ();
 fill_1 FILLER_39_275 ();
 fill_1 FILLER_39_288 ();
 fill_4 FILLER_39_309 ();
 fill_2 FILLER_39_328 ();
 fill_1 FILLER_39_356 ();
 fill_4 FILLER_39_406 ();
 fill_2 FILLER_39_431 ();
 fill_1 FILLER_39_433 ();
 fill_1 FILLER_39_447 ();
 fill_4 FILLER_39_452 ();
 fill_1 FILLER_39_456 ();
 decap_12 FILLER_39_460 ();
 fill_1 FILLER_39_472 ();
 fill_2 FILLER_39_501 ();
 fill_1 FILLER_39_503 ();
 fill_4 FILLER_39_510 ();
 fill_1 FILLER_39_514 ();
 fill_1 FILLER_39_559 ();
 fill_1 FILLER_39_594 ();
 fill_1 FILLER_39_620 ();
 fill_1 FILLER_39_642 ();
 fill_1 FILLER_39_651 ();
 fill_1 FILLER_39_671 ();
 fill_2 FILLER_39_694 ();
 fill_1 FILLER_39_721 ();
 fill_2 FILLER_39_738 ();
 fill_1 FILLER_39_803 ();
 fill_1 FILLER_39_841 ();
 fill_2 FILLER_39_868 ();
 fill_1 FILLER_39_895 ();
 fill_1 FILLER_39_903 ();
 fill_1 FILLER_39_910 ();
 fill_1 FILLER_39_951 ();
 fill_2 FILLER_39_966 ();
 fill_1 FILLER_39_1000 ();
 fill_1 FILLER_39_1024 ();
 fill_4 FILLER_39_1031 ();
 fill_2 FILLER_39_1035 ();
 fill_1 FILLER_39_1037 ();
 decap_12 FILLER_40_3 ();
 decap_12 FILLER_40_15 ();
 fill_1 FILLER_40_27 ();
 fill_1 FILLER_40_39 ();
 fill_2 FILLER_40_116 ();
 fill_1 FILLER_40_118 ();
 decap_12 FILLER_40_126 ();
 fill_2 FILLER_40_138 ();
 fill_2 FILLER_40_147 ();
 fill_2 FILLER_40_172 ();
 fill_2 FILLER_40_184 ();
 fill_2 FILLER_40_197 ();
 fill_1 FILLER_40_199 ();
 fill_1 FILLER_40_220 ();
 fill_1 FILLER_40_244 ();
 fill_2 FILLER_40_283 ();
 fill_1 FILLER_40_285 ();
 fill_1 FILLER_40_307 ();
 fill_8 FILLER_40_355 ();
 fill_1 FILLER_40_363 ();
 fill_1 FILLER_40_373 ();
 fill_1 FILLER_40_378 ();
 fill_4 FILLER_40_414 ();
 fill_2 FILLER_40_418 ();
 fill_2 FILLER_40_421 ();
 fill_1 FILLER_40_423 ();
 fill_2 FILLER_40_453 ();
 fill_2 FILLER_40_463 ();
 fill_1 FILLER_40_477 ();
 fill_4 FILLER_40_528 ();
 fill_2 FILLER_40_548 ();
 fill_1 FILLER_40_550 ();
 decap_12 FILLER_40_576 ();
 fill_8 FILLER_40_603 ();
 fill_1 FILLER_40_611 ();
 fill_2 FILLER_40_618 ();
 fill_1 FILLER_40_656 ();
 fill_1 FILLER_40_677 ();
 fill_2 FILLER_40_698 ();
 fill_1 FILLER_40_714 ();
 fill_2 FILLER_40_754 ();
 fill_2 FILLER_40_781 ();
 fill_1 FILLER_40_849 ();
 fill_1 FILLER_40_863 ();
 fill_1 FILLER_40_923 ();
 fill_2 FILLER_40_1003 ();
 fill_1 FILLER_40_1025 ();
 fill_1 FILLER_40_1035 ();
 fill_1 FILLER_40_1037 ();
 decap_12 FILLER_41_3 ();
 fill_4 FILLER_41_15 ();
 fill_1 FILLER_41_19 ();
 fill_2 FILLER_41_44 ();
 fill_2 FILLER_41_57 ();
 fill_1 FILLER_41_59 ();
 fill_2 FILLER_41_67 ();
 fill_1 FILLER_41_69 ();
 fill_8 FILLER_41_74 ();
 fill_2 FILLER_41_82 ();
 fill_2 FILLER_41_103 ();
 fill_2 FILLER_41_136 ();
 decap_12 FILLER_41_144 ();
 fill_2 FILLER_41_156 ();
 fill_2 FILLER_41_163 ();
 fill_1 FILLER_41_169 ();
 fill_2 FILLER_41_175 ();
 fill_2 FILLER_41_203 ();
 fill_2 FILLER_41_225 ();
 fill_1 FILLER_41_258 ();
 fill_2 FILLER_41_274 ();
 fill_1 FILLER_41_290 ();
 fill_4 FILLER_41_301 ();
 fill_2 FILLER_41_315 ();
 fill_1 FILLER_41_329 ();
 fill_1 FILLER_41_344 ();
 fill_2 FILLER_41_384 ();
 fill_1 FILLER_41_391 ();
 fill_1 FILLER_41_400 ();
 fill_8 FILLER_41_412 ();
 fill_1 FILLER_41_420 ();
 fill_2 FILLER_41_442 ();
 fill_1 FILLER_41_444 ();
 fill_2 FILLER_41_502 ();
 fill_2 FILLER_41_541 ();
 fill_1 FILLER_41_553 ();
 fill_1 FILLER_41_561 ();
 fill_4 FILLER_41_565 ();
 fill_2 FILLER_41_580 ();
 fill_1 FILLER_41_591 ();
 fill_2 FILLER_41_606 ();
 fill_2 FILLER_41_613 ();
 fill_1 FILLER_41_615 ();
 fill_2 FILLER_41_617 ();
 fill_1 FILLER_41_619 ();
 fill_1 FILLER_41_627 ();
 fill_2 FILLER_41_673 ();
 fill_2 FILLER_41_701 ();
 fill_1 FILLER_41_703 ();
 fill_2 FILLER_41_894 ();
 fill_2 FILLER_41_897 ();
 fill_1 FILLER_41_914 ();
 fill_1 FILLER_41_924 ();
 fill_1 FILLER_41_940 ();
 fill_1 FILLER_41_953 ();
 fill_4 FILLER_41_979 ();
 fill_2 FILLER_41_983 ();
 fill_2 FILLER_41_1006 ();
 fill_4 FILLER_41_1015 ();
 fill_2 FILLER_41_1019 ();
 fill_1 FILLER_41_1021 ();
 fill_4 FILLER_41_1031 ();
 fill_2 FILLER_41_1035 ();
 fill_1 FILLER_41_1037 ();
 decap_12 FILLER_42_3 ();
 decap_12 FILLER_42_15 ();
 fill_1 FILLER_42_27 ();
 fill_1 FILLER_42_29 ();
 fill_8 FILLER_42_46 ();
 fill_1 FILLER_42_62 ();
 fill_2 FILLER_42_82 ();
 fill_1 FILLER_42_105 ();
 fill_1 FILLER_42_123 ();
 fill_8 FILLER_42_131 ();
 fill_1 FILLER_42_139 ();
 decap_12 FILLER_42_141 ();
 decap_12 FILLER_42_153 ();
 fill_1 FILLER_42_165 ();
 fill_2 FILLER_42_181 ();
 fill_1 FILLER_42_183 ();
 fill_4 FILLER_42_197 ();
 fill_1 FILLER_42_201 ();
 fill_2 FILLER_42_217 ();
 fill_1 FILLER_42_251 ();
 fill_2 FILLER_42_268 ();
 fill_2 FILLER_42_313 ();
 fill_1 FILLER_42_363 ();
 fill_1 FILLER_42_380 ();
 fill_2 FILLER_42_412 ();
 fill_2 FILLER_42_418 ();
 fill_2 FILLER_42_441 ();
 fill_1 FILLER_42_443 ();
 fill_8 FILLER_42_458 ();
 fill_2 FILLER_42_474 ();
 fill_1 FILLER_42_508 ();
 fill_2 FILLER_42_530 ();
 fill_1 FILLER_42_549 ();
 fill_1 FILLER_42_622 ();
 fill_2 FILLER_42_671 ();
 fill_1 FILLER_42_682 ();
 fill_1 FILLER_42_688 ();
 fill_2 FILLER_42_784 ();
 fill_1 FILLER_42_797 ();
 fill_2 FILLER_42_813 ();
 fill_2 FILLER_42_842 ();
 fill_1 FILLER_42_869 ();
 fill_1 FILLER_42_923 ();
 fill_2 FILLER_42_977 ();
 fill_1 FILLER_42_979 ();
 fill_1 FILLER_42_990 ();
 fill_4 FILLER_42_1006 ();
 fill_1 FILLER_42_1010 ();
 fill_1 FILLER_42_1026 ();
 fill_1 FILLER_42_1037 ();
 decap_12 FILLER_43_3 ();
 decap_12 FILLER_43_15 ();
 fill_1 FILLER_43_27 ();
 fill_8 FILLER_43_69 ();
 fill_2 FILLER_43_77 ();
 fill_8 FILLER_43_82 ();
 fill_2 FILLER_43_90 ();
 fill_1 FILLER_43_97 ();
 fill_4 FILLER_43_136 ();
 fill_2 FILLER_43_140 ();
 fill_4 FILLER_43_149 ();
 fill_1 FILLER_43_153 ();
 fill_1 FILLER_43_167 ();
 fill_4 FILLER_43_169 ();
 fill_1 FILLER_43_173 ();
 fill_4 FILLER_43_182 ();
 fill_2 FILLER_43_186 ();
 fill_2 FILLER_43_195 ();
 fill_1 FILLER_43_197 ();
 fill_8 FILLER_43_225 ();
 fill_1 FILLER_43_233 ();
 fill_8 FILLER_43_272 ();
 fill_4 FILLER_43_288 ();
 fill_2 FILLER_43_292 ();
 fill_4 FILLER_43_300 ();
 fill_1 FILLER_43_315 ();
 fill_2 FILLER_43_326 ();
 fill_1 FILLER_43_344 ();
 fill_1 FILLER_43_384 ();
 fill_4 FILLER_43_393 ();
 fill_2 FILLER_43_397 ();
 fill_1 FILLER_43_483 ();
 fill_2 FILLER_43_502 ();
 fill_4 FILLER_43_526 ();
 fill_2 FILLER_43_534 ();
 fill_4 FILLER_43_555 ();
 fill_1 FILLER_43_559 ();
 fill_1 FILLER_43_598 ();
 fill_1 FILLER_43_651 ();
 fill_1 FILLER_43_717 ();
 fill_1 FILLER_43_727 ();
 fill_1 FILLER_43_747 ();
 fill_2 FILLER_43_841 ();
 fill_1 FILLER_43_843 ();
 fill_1 FILLER_43_856 ();
 fill_2 FILLER_43_869 ();
 fill_1 FILLER_43_891 ();
 fill_1 FILLER_43_924 ();
 fill_1 FILLER_43_943 ();
 decap_12 FILLER_44_3 ();
 decap_12 FILLER_44_15 ();
 fill_1 FILLER_44_27 ();
 fill_4 FILLER_44_51 ();
 fill_4 FILLER_44_58 ();
 fill_1 FILLER_44_78 ();
 fill_8 FILLER_44_93 ();
 decap_12 FILLER_44_119 ();
 fill_8 FILLER_44_131 ();
 fill_1 FILLER_44_139 ();
 decap_12 FILLER_44_141 ();
 fill_4 FILLER_44_153 ();
 fill_2 FILLER_44_157 ();
 fill_4 FILLER_44_162 ();
 fill_2 FILLER_44_166 ();
 fill_2 FILLER_44_220 ();
 fill_8 FILLER_44_225 ();
 fill_1 FILLER_44_233 ();
 fill_1 FILLER_44_242 ();
 fill_1 FILLER_44_251 ();
 fill_1 FILLER_44_258 ();
 fill_2 FILLER_44_296 ();
 fill_2 FILLER_44_306 ();
 fill_1 FILLER_44_317 ();
 fill_4 FILLER_44_334 ();
 fill_1 FILLER_44_338 ();
 fill_4 FILLER_44_348 ();
 fill_1 FILLER_44_352 ();
 fill_4 FILLER_44_360 ();
 fill_1 FILLER_44_365 ();
 fill_2 FILLER_44_417 ();
 fill_1 FILLER_44_419 ();
 fill_2 FILLER_44_468 ();
 fill_2 FILLER_44_494 ();
 fill_1 FILLER_44_501 ();
 fill_1 FILLER_44_515 ();
 fill_4 FILLER_44_528 ();
 decap_12 FILLER_44_575 ();
 fill_1 FILLER_44_587 ();
 fill_2 FILLER_44_589 ();
 fill_2 FILLER_44_604 ();
 fill_1 FILLER_44_668 ();
 fill_2 FILLER_44_678 ();
 fill_1 FILLER_44_725 ();
 fill_1 FILLER_44_760 ();
 fill_2 FILLER_44_813 ();
 fill_2 FILLER_44_821 ();
 fill_1 FILLER_44_867 ();
 fill_2 FILLER_44_897 ();
 fill_4 FILLER_44_920 ();
 fill_2 FILLER_44_956 ();
 fill_1 FILLER_44_958 ();
 fill_2 FILLER_44_977 ();
 fill_1 FILLER_44_979 ();
 fill_2 FILLER_44_987 ();
 fill_1 FILLER_44_1035 ();
 fill_1 FILLER_44_1037 ();
 decap_12 FILLER_45_3 ();
 fill_2 FILLER_45_15 ();
 fill_1 FILLER_45_17 ();
 fill_1 FILLER_45_26 ();
 decap_12 FILLER_45_43 ();
 fill_1 FILLER_45_55 ();
 fill_4 FILLER_45_72 ();
 fill_2 FILLER_45_76 ();
 fill_1 FILLER_45_78 ();
 fill_4 FILLER_45_86 ();
 fill_1 FILLER_45_90 ();
 fill_2 FILLER_45_106 ();
 fill_1 FILLER_45_108 ();
 fill_4 FILLER_45_117 ();
 fill_2 FILLER_45_121 ();
 fill_1 FILLER_45_123 ();
 decap_12 FILLER_45_131 ();
 fill_1 FILLER_45_143 ();
 fill_1 FILLER_45_151 ();
 fill_2 FILLER_45_159 ();
 fill_4 FILLER_45_169 ();
 fill_8 FILLER_45_177 ();
 fill_2 FILLER_45_185 ();
 fill_1 FILLER_45_187 ();
 decap_12 FILLER_45_193 ();
 fill_4 FILLER_45_205 ();
 fill_2 FILLER_45_215 ();
 fill_2 FILLER_45_245 ();
 fill_1 FILLER_45_247 ();
 fill_4 FILLER_45_256 ();
 fill_1 FILLER_45_260 ();
 fill_2 FILLER_45_322 ();
 fill_1 FILLER_45_335 ();
 fill_8 FILLER_45_362 ();
 fill_2 FILLER_45_370 ();
 decap_12 FILLER_45_380 ();
 fill_1 FILLER_45_393 ();
 fill_4 FILLER_45_443 ();
 fill_1 FILLER_45_447 ();
 fill_1 FILLER_45_458 ();
 fill_1 FILLER_45_491 ();
 fill_2 FILLER_45_501 ();
 fill_1 FILLER_45_503 ();
 fill_4 FILLER_45_513 ();
 fill_1 FILLER_45_517 ();
 fill_8 FILLER_45_529 ();
 fill_2 FILLER_45_537 ();
 decap_12 FILLER_45_561 ();
 fill_1 FILLER_45_573 ();
 fill_2 FILLER_45_594 ();
 fill_1 FILLER_45_686 ();
 fill_4 FILLER_45_710 ();
 fill_1 FILLER_45_714 ();
 fill_2 FILLER_45_735 ();
 fill_1 FILLER_45_746 ();
 fill_1 FILLER_45_783 ();
 fill_2 FILLER_45_838 ();
 fill_2 FILLER_45_841 ();
 fill_2 FILLER_45_849 ();
 fill_2 FILLER_45_857 ();
 fill_2 FILLER_45_865 ();
 fill_4 FILLER_45_921 ();
 fill_2 FILLER_45_925 ();
 fill_4 FILLER_45_936 ();
 fill_2 FILLER_45_949 ();
 fill_1 FILLER_45_951 ();
 fill_1 FILLER_45_993 ();
 fill_4 FILLER_45_1003 ();
 fill_1 FILLER_45_1007 ();
 fill_2 FILLER_45_1036 ();
 fill_2 FILLER_46_3 ();
 fill_1 FILLER_46_5 ();
 fill_1 FILLER_46_27 ();
 fill_4 FILLER_46_77 ();
 fill_2 FILLER_46_81 ();
 fill_1 FILLER_46_83 ();
 fill_8 FILLER_46_91 ();
 fill_2 FILLER_46_99 ();
 fill_4 FILLER_46_134 ();
 fill_2 FILLER_46_138 ();
 fill_8 FILLER_46_148 ();
 fill_2 FILLER_46_156 ();
 fill_4 FILLER_46_161 ();
 fill_1 FILLER_46_165 ();
 fill_2 FILLER_46_173 ();
 fill_4 FILLER_46_182 ();
 fill_1 FILLER_46_186 ();
 fill_2 FILLER_46_194 ();
 fill_1 FILLER_46_215 ();
 decap_12 FILLER_46_223 ();
 decap_12 FILLER_46_235 ();
 fill_4 FILLER_46_247 ();
 fill_1 FILLER_46_251 ();
 decap_12 FILLER_46_253 ();
 decap_12 FILLER_46_265 ();
 fill_4 FILLER_46_277 ();
 fill_2 FILLER_46_281 ();
 fill_1 FILLER_46_294 ();
 fill_1 FILLER_46_298 ();
 fill_1 FILLER_46_307 ();
 fill_8 FILLER_46_309 ();
 fill_2 FILLER_46_317 ();
 fill_2 FILLER_46_331 ();
 fill_2 FILLER_46_352 ();
 fill_1 FILLER_46_354 ();
 fill_1 FILLER_46_363 ();
 fill_2 FILLER_46_372 ();
 fill_1 FILLER_46_374 ();
 fill_1 FILLER_46_382 ();
 fill_1 FILLER_46_410 ();
 fill_4 FILLER_46_416 ();
 fill_2 FILLER_46_444 ();
 fill_2 FILLER_46_474 ();
 fill_1 FILLER_46_485 ();
 fill_2 FILLER_46_507 ();
 fill_1 FILLER_46_509 ();
 fill_1 FILLER_46_531 ();
 fill_4 FILLER_46_538 ();
 fill_2 FILLER_46_542 ();
 fill_4 FILLER_46_554 ();
 fill_1 FILLER_46_558 ();
 fill_2 FILLER_46_562 ();
 fill_1 FILLER_46_564 ();
 fill_4 FILLER_46_578 ();
 fill_2 FILLER_46_582 ();
 fill_1 FILLER_46_587 ();
 fill_2 FILLER_46_594 ();
 fill_2 FILLER_46_611 ();
 fill_2 FILLER_46_684 ();
 fill_1 FILLER_46_686 ();
 fill_1 FILLER_46_705 ();
 fill_2 FILLER_46_754 ();
 fill_2 FILLER_46_842 ();
 fill_2 FILLER_46_853 ();
 fill_1 FILLER_46_855 ();
 fill_2 FILLER_46_905 ();
 fill_4 FILLER_46_919 ();
 fill_1 FILLER_46_923 ();
 fill_2 FILLER_46_978 ();
 fill_1 FILLER_46_1037 ();
 fill_4 FILLER_47_3 ();
 fill_2 FILLER_47_7 ();
 fill_1 FILLER_47_9 ();
 fill_4 FILLER_47_32 ();
 fill_1 FILLER_47_36 ();
 fill_4 FILLER_47_44 ();
 fill_1 FILLER_47_48 ();
 fill_2 FILLER_47_57 ();
 fill_1 FILLER_47_59 ();
 fill_2 FILLER_47_101 ();
 fill_1 FILLER_47_111 ();
 fill_2 FILLER_47_118 ();
 fill_1 FILLER_47_120 ();
 decap_12 FILLER_47_128 ();
 fill_8 FILLER_47_140 ();
 fill_2 FILLER_47_148 ();
 fill_8 FILLER_47_157 ();
 fill_2 FILLER_47_165 ();
 fill_1 FILLER_47_167 ();
 decap_12 FILLER_47_182 ();
 decap_12 FILLER_47_194 ();
 fill_4 FILLER_47_206 ();
 fill_1 FILLER_47_210 ();
 fill_4 FILLER_47_218 ();
 fill_2 FILLER_47_222 ();
 decap_12 FILLER_47_225 ();
 fill_1 FILLER_47_237 ();
 decap_12 FILLER_47_245 ();
 fill_2 FILLER_47_257 ();
 fill_1 FILLER_47_259 ();
 decap_12 FILLER_47_267 ();
 fill_1 FILLER_47_279 ();
 fill_1 FILLER_47_307 ();
 fill_2 FILLER_47_316 ();
 fill_2 FILLER_47_334 ();
 fill_4 FILLER_47_345 ();
 fill_2 FILLER_47_349 ();
 fill_2 FILLER_47_377 ();
 fill_1 FILLER_47_379 ();
 fill_1 FILLER_47_391 ();
 fill_2 FILLER_47_393 ();
 fill_1 FILLER_47_395 ();
 fill_2 FILLER_47_422 ();
 fill_1 FILLER_47_424 ();
 decap_12 FILLER_47_434 ();
 fill_2 FILLER_47_446 ();
 fill_1 FILLER_47_484 ();
 fill_2 FILLER_47_501 ();
 fill_1 FILLER_47_503 ();
 fill_1 FILLER_47_524 ();
 fill_2 FILLER_47_558 ();
 fill_2 FILLER_47_577 ();
 fill_2 FILLER_47_679 ();
 fill_1 FILLER_47_681 ();
 fill_2 FILLER_47_700 ();
 fill_1 FILLER_47_702 ();
 fill_1 FILLER_47_723 ();
 fill_2 FILLER_47_744 ();
 fill_2 FILLER_47_791 ();
 fill_1 FILLER_47_813 ();
 fill_2 FILLER_47_835 ();
 fill_1 FILLER_47_932 ();
 fill_1 FILLER_47_951 ();
 fill_2 FILLER_47_962 ();
 fill_2 FILLER_47_990 ();
 fill_2 FILLER_47_1002 ();
 fill_1 FILLER_47_1004 ();
 fill_2 FILLER_47_1009 ();
 fill_1 FILLER_48_27 ();
 fill_4 FILLER_48_52 ();
 fill_2 FILLER_48_56 ();
 fill_1 FILLER_48_66 ();
 fill_4 FILLER_48_128 ();
 fill_1 FILLER_48_132 ();
 fill_1 FILLER_48_141 ();
 fill_4 FILLER_48_149 ();
 fill_1 FILLER_48_153 ();
 fill_4 FILLER_48_161 ();
 decap_12 FILLER_48_168 ();
 fill_2 FILLER_48_180 ();
 fill_1 FILLER_48_182 ();
 fill_4 FILLER_48_190 ();
 fill_2 FILLER_48_194 ();
 fill_8 FILLER_48_197 ();
 fill_2 FILLER_48_205 ();
 fill_8 FILLER_48_214 ();
 fill_1 FILLER_48_222 ();
 decap_12 FILLER_48_230 ();
 fill_8 FILLER_48_242 ();
 fill_2 FILLER_48_250 ();
 decap_12 FILLER_48_253 ();
 fill_4 FILLER_48_265 ();
 fill_2 FILLER_48_269 ();
 fill_8 FILLER_48_278 ();
 fill_1 FILLER_48_286 ();
 fill_1 FILLER_48_294 ();
 fill_2 FILLER_48_306 ();
 fill_8 FILLER_48_330 ();
 fill_1 FILLER_48_338 ();
 fill_2 FILLER_48_354 ();
 fill_2 FILLER_48_365 ();
 fill_1 FILLER_48_367 ();
 fill_1 FILLER_48_375 ();
 fill_4 FILLER_48_380 ();
 fill_2 FILLER_48_384 ();
 fill_1 FILLER_48_386 ();
 fill_8 FILLER_48_394 ();
 fill_4 FILLER_48_406 ();
 fill_1 FILLER_48_410 ();
 fill_4 FILLER_48_414 ();
 fill_2 FILLER_48_418 ();
 fill_4 FILLER_48_445 ();
 fill_2 FILLER_48_449 ();
 fill_8 FILLER_48_477 ();
 fill_2 FILLER_48_485 ();
 fill_1 FILLER_48_487 ();
 fill_2 FILLER_48_499 ();
 fill_1 FILLER_48_505 ();
 fill_4 FILLER_48_510 ();
 fill_2 FILLER_48_514 ();
 fill_2 FILLER_48_533 ();
 fill_1 FILLER_48_543 ();
 decap_12 FILLER_48_559 ();
 fill_4 FILLER_48_571 ();
 fill_2 FILLER_48_595 ();
 fill_1 FILLER_48_597 ();
 fill_1 FILLER_48_634 ();
 fill_1 FILLER_48_643 ();
 fill_1 FILLER_48_710 ();
 fill_1 FILLER_48_769 ();
 fill_2 FILLER_48_839 ();
 fill_2 FILLER_48_865 ();
 fill_1 FILLER_48_867 ();
 fill_8 FILLER_48_869 ();
 fill_2 FILLER_48_877 ();
 fill_1 FILLER_48_879 ();
 fill_1 FILLER_48_923 ();
 fill_1 FILLER_48_925 ();
 fill_1 FILLER_48_979 ();
 fill_2 FILLER_48_999 ();
 fill_1 FILLER_48_1013 ();
 fill_2 FILLER_48_1034 ();
 fill_1 FILLER_48_1037 ();
 fill_8 FILLER_49_3 ();
 fill_2 FILLER_49_30 ();
 fill_2 FILLER_49_39 ();
 fill_1 FILLER_49_41 ();
 fill_2 FILLER_49_46 ();
 fill_1 FILLER_49_48 ();
 fill_4 FILLER_49_83 ();
 fill_2 FILLER_49_87 ();
 fill_2 FILLER_49_110 ();
 decap_12 FILLER_49_117 ();
 fill_1 FILLER_49_129 ();
 decap_12 FILLER_49_133 ();
 decap_12 FILLER_49_145 ();
 fill_4 FILLER_49_157 ();
 fill_1 FILLER_49_169 ();
 fill_4 FILLER_49_177 ();
 fill_1 FILLER_49_191 ();
 fill_8 FILLER_49_207 ();
 fill_2 FILLER_49_215 ();
 fill_4 FILLER_49_229 ();
 fill_2 FILLER_49_233 ();
 fill_1 FILLER_49_235 ();
 fill_4 FILLER_49_243 ();
 fill_2 FILLER_49_247 ();
 fill_2 FILLER_49_256 ();
 fill_1 FILLER_49_258 ();
 fill_4 FILLER_49_266 ();
 fill_1 FILLER_49_270 ();
 fill_4 FILLER_49_275 ();
 fill_1 FILLER_49_279 ();
 decap_12 FILLER_49_281 ();
 decap_12 FILLER_49_293 ();
 decap_12 FILLER_49_305 ();
 fill_4 FILLER_49_324 ();
 fill_1 FILLER_49_328 ();
 fill_1 FILLER_49_345 ();
 fill_1 FILLER_49_355 ();
 fill_2 FILLER_49_420 ();
 fill_4 FILLER_49_472 ();
 fill_4 FILLER_49_483 ();
 fill_2 FILLER_49_494 ();
 fill_1 FILLER_49_556 ();
 fill_4 FILLER_49_572 ();
 fill_2 FILLER_49_576 ();
 fill_2 FILLER_49_586 ();
 fill_1 FILLER_49_588 ();
 fill_4 FILLER_49_596 ();
 fill_1 FILLER_49_617 ();
 fill_2 FILLER_49_679 ();
 fill_4 FILLER_49_687 ();
 fill_1 FILLER_49_697 ();
 fill_4 FILLER_49_748 ();
 fill_1 FILLER_49_756 ();
 fill_2 FILLER_49_779 ();
 fill_2 FILLER_49_812 ();
 fill_2 FILLER_49_844 ();
 fill_2 FILLER_49_849 ();
 fill_2 FILLER_49_871 ();
 fill_1 FILLER_49_873 ();
 fill_2 FILLER_49_894 ();
 fill_1 FILLER_49_910 ();
 fill_4 FILLER_49_931 ();
 fill_1 FILLER_49_935 ();
 fill_8 FILLER_49_942 ();
 fill_2 FILLER_49_950 ();
 fill_1 FILLER_49_979 ();
 fill_4 FILLER_49_1003 ();
 fill_1 FILLER_49_1007 ();
 fill_4 FILLER_49_1018 ();
 fill_1 FILLER_49_1022 ();
 fill_1 FILLER_50_19 ();
 fill_1 FILLER_50_27 ();
 fill_4 FILLER_50_33 ();
 fill_1 FILLER_50_45 ();
 fill_4 FILLER_50_50 ();
 fill_2 FILLER_50_54 ();
 fill_1 FILLER_50_56 ();
 fill_2 FILLER_50_72 ();
 fill_1 FILLER_50_74 ();
 fill_2 FILLER_50_82 ();
 fill_2 FILLER_50_89 ();
 fill_2 FILLER_50_108 ();
 fill_2 FILLER_50_126 ();
 fill_2 FILLER_50_137 ();
 fill_1 FILLER_50_139 ();
 fill_4 FILLER_50_148 ();
 decap_12 FILLER_50_168 ();
 decap_12 FILLER_50_180 ();
 fill_4 FILLER_50_192 ();
 decap_12 FILLER_50_197 ();
 fill_2 FILLER_50_209 ();
 decap_12 FILLER_50_218 ();
 fill_4 FILLER_50_230 ();
 fill_8 FILLER_50_242 ();
 fill_2 FILLER_50_250 ();
 decap_12 FILLER_50_253 ();
 fill_4 FILLER_50_265 ();
 fill_2 FILLER_50_269 ();
 fill_1 FILLER_50_271 ();
 fill_2 FILLER_50_286 ();
 fill_1 FILLER_50_288 ();
 fill_2 FILLER_50_361 ();
 fill_1 FILLER_50_363 ();
 fill_8 FILLER_50_365 ();
 fill_1 FILLER_50_373 ();
 fill_8 FILLER_50_378 ();
 fill_2 FILLER_50_386 ();
 fill_8 FILLER_50_393 ();
 fill_2 FILLER_50_401 ();
 fill_8 FILLER_50_489 ();
 fill_1 FILLER_50_497 ();
 fill_4 FILLER_50_528 ();
 fill_2 FILLER_50_541 ();
 fill_1 FILLER_50_543 ();
 fill_4 FILLER_50_589 ();
 fill_1 FILLER_50_622 ();
 fill_1 FILLER_50_657 ();
 fill_2 FILLER_50_710 ();
 fill_1 FILLER_50_712 ();
 fill_4 FILLER_50_735 ();
 fill_1 FILLER_50_739 ();
 fill_1 FILLER_50_755 ();
 fill_8 FILLER_50_819 ();
 fill_2 FILLER_50_836 ();
 fill_1 FILLER_50_838 ();
 fill_2 FILLER_50_866 ();
 fill_2 FILLER_50_869 ();
 fill_1 FILLER_50_892 ();
 fill_1 FILLER_50_896 ();
 fill_1 FILLER_50_906 ();
 fill_2 FILLER_50_922 ();
 fill_2 FILLER_50_928 ();
 fill_4 FILLER_50_936 ();
 fill_2 FILLER_50_969 ();
 fill_1 FILLER_50_981 ();
 fill_2 FILLER_50_985 ();
 fill_1 FILLER_50_987 ();
 fill_2 FILLER_50_1003 ();
 fill_1 FILLER_50_1005 ();
 fill_2 FILLER_50_1015 ();
 fill_1 FILLER_50_1017 ();
 fill_1 FILLER_50_1037 ();
 fill_4 FILLER_51_3 ();
 fill_1 FILLER_51_7 ();
 fill_1 FILLER_51_18 ();
 fill_2 FILLER_51_26 ();
 fill_1 FILLER_51_61 ();
 fill_1 FILLER_51_71 ();
 fill_1 FILLER_51_85 ();
 fill_4 FILLER_51_93 ();
 fill_2 FILLER_51_97 ();
 fill_4 FILLER_51_105 ();
 fill_2 FILLER_51_109 ();
 fill_1 FILLER_51_111 ();
 fill_2 FILLER_51_116 ();
 fill_4 FILLER_51_156 ();
 fill_1 FILLER_51_167 ();
 fill_2 FILLER_51_169 ();
 fill_1 FILLER_51_171 ();
 fill_2 FILLER_51_180 ();
 fill_1 FILLER_51_182 ();
 fill_1 FILLER_51_190 ();
 decap_12 FILLER_51_206 ();
 fill_4 FILLER_51_218 ();
 fill_2 FILLER_51_222 ();
 fill_4 FILLER_51_225 ();
 fill_1 FILLER_51_229 ();
 decap_12 FILLER_51_235 ();
 fill_8 FILLER_51_247 ();
 fill_2 FILLER_51_255 ();
 fill_1 FILLER_51_257 ();
 decap_12 FILLER_51_265 ();
 fill_2 FILLER_51_277 ();
 fill_1 FILLER_51_279 ();
 decap_12 FILLER_51_281 ();
 fill_4 FILLER_51_293 ();
 fill_8 FILLER_51_305 ();
 fill_1 FILLER_51_320 ();
 fill_8 FILLER_51_325 ();
 fill_2 FILLER_51_333 ();
 fill_1 FILLER_51_335 ();
 fill_4 FILLER_51_337 ();
 fill_2 FILLER_51_341 ();
 fill_4 FILLER_51_351 ();
 fill_4 FILLER_51_378 ();
 fill_2 FILLER_51_382 ();
 fill_1 FILLER_51_391 ();
 fill_8 FILLER_51_449 ();
 decap_12 FILLER_51_466 ();
 decap_12 FILLER_51_492 ();
 fill_1 FILLER_51_513 ();
 fill_4 FILLER_51_561 ();
 fill_1 FILLER_51_565 ();
 fill_1 FILLER_51_671 ();
 fill_2 FILLER_51_726 ();
 fill_2 FILLER_51_742 ();
 fill_1 FILLER_51_744 ();
 fill_1 FILLER_51_783 ();
 fill_1 FILLER_51_785 ();
 fill_1 FILLER_51_807 ();
 fill_2 FILLER_51_811 ();
 fill_1 FILLER_51_833 ();
 fill_4 FILLER_51_850 ();
 fill_1 FILLER_51_854 ();
 fill_2 FILLER_51_887 ();
 fill_1 FILLER_51_889 ();
 fill_1 FILLER_51_906 ();
 fill_2 FILLER_51_950 ();
 fill_1 FILLER_51_953 ();
 fill_2 FILLER_51_986 ();
 fill_4 FILLER_51_1009 ();
 fill_1 FILLER_51_1013 ();
 fill_1 FILLER_51_1037 ();
 fill_2 FILLER_52_19 ();
 fill_1 FILLER_52_21 ();
 fill_2 FILLER_52_26 ();
 decap_12 FILLER_52_29 ();
 fill_2 FILLER_52_41 ();
 fill_1 FILLER_52_77 ();
 fill_1 FILLER_52_83 ();
 fill_2 FILLER_52_85 ();
 fill_1 FILLER_52_87 ();
 fill_2 FILLER_52_107 ();
 fill_4 FILLER_52_113 ();
 fill_2 FILLER_52_117 ();
 decap_12 FILLER_52_128 ();
 fill_4 FILLER_52_141 ();
 fill_1 FILLER_52_145 ();
 fill_2 FILLER_52_150 ();
 fill_1 FILLER_52_152 ();
 fill_2 FILLER_52_175 ();
 decap_12 FILLER_52_184 ();
 fill_2 FILLER_52_197 ();
 fill_1 FILLER_52_206 ();
 fill_4 FILLER_52_224 ();
 fill_2 FILLER_52_228 ();
 fill_4 FILLER_52_239 ();
 fill_1 FILLER_52_243 ();
 fill_1 FILLER_52_251 ();
 decap_12 FILLER_52_273 ();
 fill_4 FILLER_52_285 ();
 fill_2 FILLER_52_309 ();
 fill_1 FILLER_52_311 ();
 fill_1 FILLER_52_353 ();
 fill_2 FILLER_52_362 ();
 fill_2 FILLER_52_365 ();
 fill_1 FILLER_52_378 ();
 fill_1 FILLER_52_419 ();
 fill_1 FILLER_52_421 ();
 fill_2 FILLER_52_431 ();
 fill_4 FILLER_52_472 ();
 decap_12 FILLER_52_477 ();
 fill_1 FILLER_52_489 ();
 fill_1 FILLER_52_531 ();
 fill_2 FILLER_52_559 ();
 fill_1 FILLER_52_587 ();
 fill_1 FILLER_52_755 ();
 fill_1 FILLER_52_811 ();
 fill_1 FILLER_52_834 ();
 fill_2 FILLER_52_855 ();
 fill_2 FILLER_52_866 ();
 fill_4 FILLER_52_869 ();
 fill_2 FILLER_52_873 ();
 fill_1 FILLER_52_875 ();
 fill_4 FILLER_52_916 ();
 fill_1 FILLER_52_920 ();
 fill_1 FILLER_52_955 ();
 fill_1 FILLER_52_1005 ();
 fill_2 FILLER_52_1033 ();
 fill_1 FILLER_52_1035 ();
 fill_1 FILLER_52_1037 ();
 fill_1 FILLER_53_3 ();
 fill_2 FILLER_53_54 ();
 fill_8 FILLER_53_57 ();
 fill_2 FILLER_53_65 ();
 decap_12 FILLER_53_122 ();
 decap_12 FILLER_53_134 ();
 fill_8 FILLER_53_151 ();
 fill_2 FILLER_53_166 ();
 decap_12 FILLER_53_169 ();
 fill_8 FILLER_53_181 ();
 fill_1 FILLER_53_189 ();
 decap_12 FILLER_53_196 ();
 decap_12 FILLER_53_208 ();
 fill_4 FILLER_53_220 ();
 fill_1 FILLER_53_225 ();
 decap_12 FILLER_53_234 ();
 fill_8 FILLER_53_246 ();
 fill_1 FILLER_53_254 ();
 fill_8 FILLER_53_267 ();
 fill_1 FILLER_53_275 ();
 fill_1 FILLER_53_326 ();
 fill_2 FILLER_53_333 ();
 fill_1 FILLER_53_335 ();
 fill_4 FILLER_53_337 ();
 fill_1 FILLER_53_341 ();
 fill_4 FILLER_53_357 ();
 fill_1 FILLER_53_361 ();
 fill_2 FILLER_53_369 ();
 fill_4 FILLER_53_378 ();
 fill_1 FILLER_53_382 ();
 fill_2 FILLER_53_390 ();
 fill_1 FILLER_53_396 ();
 fill_1 FILLER_53_411 ();
 fill_2 FILLER_53_428 ();
 fill_4 FILLER_53_449 ();
 fill_2 FILLER_53_453 ();
 decap_12 FILLER_53_473 ();
 fill_1 FILLER_53_496 ();
 fill_2 FILLER_53_513 ();
 fill_1 FILLER_53_531 ();
 fill_2 FILLER_53_541 ();
 fill_2 FILLER_53_585 ();
 fill_1 FILLER_53_595 ();
 fill_1 FILLER_53_606 ();
 fill_1 FILLER_53_646 ();
 fill_2 FILLER_53_655 ();
 fill_1 FILLER_53_657 ();
 fill_8 FILLER_53_673 ();
 fill_2 FILLER_53_681 ();
 fill_2 FILLER_53_701 ();
 fill_1 FILLER_53_763 ();
 fill_1 FILLER_53_791 ();
 fill_2 FILLER_53_903 ();
 fill_2 FILLER_53_924 ();
 fill_4 FILLER_53_962 ();
 fill_2 FILLER_53_966 ();
 fill_8 FILLER_53_991 ();
 fill_2 FILLER_53_1012 ();
 fill_1 FILLER_53_1037 ();
 fill_8 FILLER_54_3 ();
 fill_1 FILLER_54_15 ();
 fill_4 FILLER_54_23 ();
 fill_1 FILLER_54_27 ();
 fill_8 FILLER_54_29 ();
 fill_2 FILLER_54_37 ();
 fill_1 FILLER_54_39 ();
 fill_4 FILLER_54_60 ();
 fill_2 FILLER_54_64 ();
 fill_1 FILLER_54_71 ();
 fill_4 FILLER_54_80 ();
 fill_4 FILLER_54_90 ();
 fill_2 FILLER_54_94 ();
 fill_1 FILLER_54_96 ();
 fill_1 FILLER_54_102 ();
 fill_4 FILLER_54_124 ();
 fill_1 FILLER_54_128 ();
 fill_2 FILLER_54_137 ();
 fill_1 FILLER_54_139 ();
 fill_8 FILLER_54_160 ();
 fill_8 FILLER_54_173 ();
 fill_8 FILLER_54_185 ();
 fill_2 FILLER_54_193 ();
 fill_1 FILLER_54_195 ();
 fill_2 FILLER_54_211 ();
 decap_12 FILLER_54_217 ();
 fill_2 FILLER_54_229 ();
 fill_1 FILLER_54_231 ();
 fill_4 FILLER_54_239 ();
 fill_4 FILLER_54_248 ();
 fill_2 FILLER_54_260 ();
 fill_1 FILLER_54_262 ();
 fill_2 FILLER_54_284 ();
 fill_2 FILLER_54_302 ();
 fill_2 FILLER_54_317 ();
 fill_8 FILLER_54_327 ();
 fill_2 FILLER_54_335 ();
 fill_1 FILLER_54_337 ();
 fill_4 FILLER_54_346 ();
 fill_1 FILLER_54_350 ();
 fill_2 FILLER_54_362 ();
 fill_1 FILLER_54_365 ();
 fill_2 FILLER_54_417 ();
 fill_1 FILLER_54_419 ();
 fill_1 FILLER_54_430 ();
 fill_2 FILLER_54_440 ();
 fill_1 FILLER_54_442 ();
 fill_4 FILLER_54_452 ();
 fill_1 FILLER_54_456 ();
 fill_2 FILLER_54_466 ();
 fill_1 FILLER_54_477 ();
 fill_1 FILLER_54_487 ();
 fill_4 FILLER_54_493 ();
 fill_2 FILLER_54_533 ();
 fill_2 FILLER_54_546 ();
 fill_1 FILLER_54_596 ();
 fill_1 FILLER_54_630 ();
 fill_2 FILLER_54_677 ();
 fill_1 FILLER_54_679 ();
 fill_2 FILLER_54_689 ();
 fill_1 FILLER_54_775 ();
 fill_1 FILLER_54_789 ();
 fill_1 FILLER_54_867 ();
 fill_1 FILLER_54_893 ();
 fill_1 FILLER_54_903 ();
 fill_4 FILLER_54_929 ();
 fill_2 FILLER_54_977 ();
 fill_1 FILLER_54_979 ();
 fill_1 FILLER_54_990 ();
 decap_12 FILLER_54_1021 ();
 fill_1 FILLER_54_1037 ();
 decap_12 FILLER_55_24 ();
 fill_2 FILLER_55_47 ();
 fill_2 FILLER_55_53 ();
 fill_1 FILLER_55_55 ();
 fill_2 FILLER_55_57 ();
 fill_4 FILLER_55_77 ();
 fill_2 FILLER_55_96 ();
 fill_1 FILLER_55_111 ();
 fill_4 FILLER_55_126 ();
 fill_2 FILLER_55_130 ();
 decap_12 FILLER_55_139 ();
 fill_2 FILLER_55_151 ();
 fill_2 FILLER_55_165 ();
 fill_1 FILLER_55_167 ();
 fill_8 FILLER_55_176 ();
 fill_2 FILLER_55_184 ();
 decap_12 FILLER_55_193 ();
 fill_4 FILLER_55_205 ();
 fill_8 FILLER_55_216 ();
 decap_12 FILLER_55_232 ();
 fill_4 FILLER_55_244 ();
 fill_1 FILLER_55_248 ();
 fill_1 FILLER_55_256 ();
 fill_2 FILLER_55_264 ();
 fill_1 FILLER_55_266 ();
 fill_4 FILLER_55_274 ();
 fill_2 FILLER_55_278 ();
 fill_4 FILLER_55_294 ();
 fill_1 FILLER_55_328 ();
 fill_2 FILLER_55_367 ();
 fill_2 FILLER_55_380 ();
 fill_1 FILLER_55_382 ();
 fill_2 FILLER_55_390 ();
 fill_1 FILLER_55_408 ();
 fill_1 FILLER_55_437 ();
 fill_1 FILLER_55_474 ();
 fill_8 FILLER_55_487 ();
 fill_1 FILLER_55_495 ();
 fill_1 FILLER_55_514 ();
 fill_2 FILLER_55_520 ();
 fill_2 FILLER_55_527 ();
 fill_4 FILLER_55_534 ();
 fill_2 FILLER_55_546 ();
 fill_4 FILLER_55_556 ();
 fill_2 FILLER_55_569 ();
 fill_2 FILLER_55_608 ();
 fill_2 FILLER_55_664 ();
 fill_1 FILLER_55_696 ();
 fill_1 FILLER_55_727 ();
 fill_2 FILLER_55_766 ();
 fill_1 FILLER_55_783 ();
 fill_1 FILLER_55_805 ();
 fill_1 FILLER_55_835 ();
 fill_2 FILLER_55_871 ();
 fill_2 FILLER_55_894 ();
 fill_1 FILLER_55_937 ();
 fill_4 FILLER_55_947 ();
 fill_1 FILLER_55_951 ();
 fill_2 FILLER_55_956 ();
 fill_1 FILLER_55_958 ();
 fill_2 FILLER_55_991 ();
 fill_4 FILLER_55_1009 ();
 fill_2 FILLER_55_1013 ();
 fill_1 FILLER_55_1015 ();
 fill_8 FILLER_55_1028 ();
 fill_2 FILLER_55_1036 ();
 fill_4 FILLER_56_3 ();
 fill_2 FILLER_56_7 ();
 fill_2 FILLER_56_29 ();
 fill_8 FILLER_56_50 ();
 fill_1 FILLER_56_58 ();
 fill_8 FILLER_56_76 ();
 fill_2 FILLER_56_104 ();
 fill_1 FILLER_56_125 ();
 fill_4 FILLER_56_133 ();
 fill_2 FILLER_56_137 ();
 fill_1 FILLER_56_139 ();
 fill_2 FILLER_56_141 ();
 fill_1 FILLER_56_143 ();
 fill_1 FILLER_56_148 ();
 fill_4 FILLER_56_156 ();
 fill_4 FILLER_56_167 ();
 fill_1 FILLER_56_171 ();
 fill_8 FILLER_56_186 ();
 fill_2 FILLER_56_194 ();
 fill_2 FILLER_56_197 ();
 fill_1 FILLER_56_199 ();
 decap_12 FILLER_56_205 ();
 fill_1 FILLER_56_217 ();
 fill_8 FILLER_56_224 ();
 fill_2 FILLER_56_232 ();
 fill_4 FILLER_56_241 ();
 fill_2 FILLER_56_245 ();
 fill_2 FILLER_56_250 ();
 fill_2 FILLER_56_253 ();
 fill_2 FILLER_56_269 ();
 fill_1 FILLER_56_271 ();
 fill_1 FILLER_56_286 ();
 fill_8 FILLER_56_299 ();
 fill_1 FILLER_56_307 ();
 fill_4 FILLER_56_309 ();
 fill_2 FILLER_56_313 ();
 fill_2 FILLER_56_325 ();
 fill_1 FILLER_56_327 ();
 fill_4 FILLER_56_334 ();
 fill_2 FILLER_56_338 ();
 fill_1 FILLER_56_340 ();
 fill_2 FILLER_56_348 ();
 fill_1 FILLER_56_350 ();
 fill_8 FILLER_56_356 ();
 fill_1 FILLER_56_365 ();
 fill_4 FILLER_56_374 ();
 fill_2 FILLER_56_378 ();
 decap_12 FILLER_56_408 ();
 fill_8 FILLER_56_421 ();
 fill_2 FILLER_56_429 ();
 fill_4 FILLER_56_445 ();
 fill_2 FILLER_56_449 ();
 fill_1 FILLER_56_451 ();
 fill_2 FILLER_56_461 ();
 fill_2 FILLER_56_480 ();
 fill_1 FILLER_56_482 ();
 fill_2 FILLER_56_498 ();
 fill_1 FILLER_56_508 ();
 fill_1 FILLER_56_521 ();
 fill_2 FILLER_56_529 ();
 fill_1 FILLER_56_531 ();
 fill_2 FILLER_56_533 ();
 fill_1 FILLER_56_535 ();
 fill_4 FILLER_56_547 ();
 fill_1 FILLER_56_564 ();
 fill_2 FILLER_56_586 ();
 fill_2 FILLER_56_642 ();
 fill_1 FILLER_56_674 ();
 fill_2 FILLER_56_698 ();
 fill_2 FILLER_56_713 ();
 fill_1 FILLER_56_715 ();
 fill_1 FILLER_56_769 ();
 fill_1 FILLER_56_805 ();
 fill_1 FILLER_56_855 ();
 fill_1 FILLER_56_960 ();
 fill_1 FILLER_56_981 ();
 fill_1 FILLER_56_1037 ();
 fill_2 FILLER_57_3 ();
 fill_1 FILLER_57_40 ();
 fill_4 FILLER_57_44 ();
 fill_1 FILLER_57_48 ();
 fill_2 FILLER_57_53 ();
 fill_1 FILLER_57_55 ();
 fill_2 FILLER_57_73 ();
 fill_1 FILLER_57_75 ();
 fill_2 FILLER_57_81 ();
 fill_1 FILLER_57_90 ();
 fill_2 FILLER_57_109 ();
 fill_1 FILLER_57_111 ();
 fill_8 FILLER_57_121 ();
 fill_2 FILLER_57_129 ();
 decap_12 FILLER_57_138 ();
 fill_1 FILLER_57_150 ();
 fill_2 FILLER_57_166 ();
 fill_1 FILLER_57_169 ();
 fill_4 FILLER_57_183 ();
 fill_4 FILLER_57_194 ();
 fill_4 FILLER_57_220 ();
 fill_4 FILLER_57_225 ();
 fill_2 FILLER_57_240 ();
 fill_1 FILLER_57_273 ();
 fill_2 FILLER_57_294 ();
 fill_2 FILLER_57_326 ();
 fill_1 FILLER_57_362 ();
 fill_4 FILLER_57_387 ();
 fill_1 FILLER_57_391 ();
 fill_2 FILLER_57_393 ();
 fill_1 FILLER_57_395 ();
 fill_4 FILLER_57_444 ();
 fill_1 FILLER_57_468 ();
 fill_8 FILLER_57_481 ();
 fill_2 FILLER_57_489 ();
 fill_4 FILLER_57_500 ();
 fill_1 FILLER_57_510 ();
 fill_4 FILLER_57_520 ();
 fill_1 FILLER_57_524 ();
 fill_8 FILLER_57_532 ();
 fill_2 FILLER_57_558 ();
 fill_1 FILLER_57_591 ();
 fill_1 FILLER_57_612 ();
 fill_1 FILLER_57_637 ();
 fill_2 FILLER_57_698 ();
 fill_4 FILLER_57_723 ();
 fill_1 FILLER_57_727 ();
 fill_4 FILLER_57_757 ();
 fill_1 FILLER_57_761 ();
 fill_2 FILLER_57_782 ();
 fill_2 FILLER_57_808 ();
 fill_1 FILLER_57_833 ();
 fill_2 FILLER_57_894 ();
 fill_1 FILLER_57_936 ();
 fill_4 FILLER_57_1017 ();
 fill_1 FILLER_57_1021 ();
 fill_4 FILLER_57_1031 ();
 fill_2 FILLER_57_1035 ();
 fill_1 FILLER_57_1037 ();
 fill_2 FILLER_58_19 ();
 fill_1 FILLER_58_50 ();
 fill_1 FILLER_58_65 ();
 fill_1 FILLER_58_83 ();
 fill_1 FILLER_58_112 ();
 fill_8 FILLER_58_131 ();
 fill_1 FILLER_58_139 ();
 fill_4 FILLER_58_141 ();
 fill_1 FILLER_58_145 ();
 decap_12 FILLER_58_154 ();
 fill_2 FILLER_58_166 ();
 fill_1 FILLER_58_168 ();
 fill_2 FILLER_58_181 ();
 fill_4 FILLER_58_190 ();
 fill_2 FILLER_58_194 ();
 fill_4 FILLER_58_197 ();
 fill_2 FILLER_58_201 ();
 fill_2 FILLER_58_212 ();
 fill_2 FILLER_58_228 ();
 fill_1 FILLER_58_230 ();
 fill_4 FILLER_58_240 ();
 fill_2 FILLER_58_249 ();
 fill_1 FILLER_58_251 ();
 fill_8 FILLER_58_253 ();
 fill_1 FILLER_58_269 ();
 fill_1 FILLER_58_273 ();
 fill_8 FILLER_58_299 ();
 fill_1 FILLER_58_307 ();
 fill_4 FILLER_58_309 ();
 fill_1 FILLER_58_313 ();
 fill_4 FILLER_58_337 ();
 fill_2 FILLER_58_349 ();
 fill_4 FILLER_58_358 ();
 fill_2 FILLER_58_362 ();
 fill_1 FILLER_58_365 ();
 fill_1 FILLER_58_376 ();
 fill_4 FILLER_58_389 ();
 fill_1 FILLER_58_410 ();
 fill_4 FILLER_58_446 ();
 fill_2 FILLER_58_459 ();
 fill_1 FILLER_58_461 ();
 fill_1 FILLER_58_480 ();
 fill_4 FILLER_58_488 ();
 fill_2 FILLER_58_492 ();
 fill_4 FILLER_58_500 ();
 fill_2 FILLER_58_504 ();
 fill_1 FILLER_58_506 ();
 fill_8 FILLER_58_511 ();
 fill_2 FILLER_58_519 ();
 fill_4 FILLER_58_528 ();
 decap_12 FILLER_58_606 ();
 fill_1 FILLER_58_618 ();
 fill_2 FILLER_58_629 ();
 fill_1 FILLER_58_645 ();
 fill_2 FILLER_58_697 ();
 fill_1 FILLER_58_699 ();
 fill_4 FILLER_58_709 ();
 fill_2 FILLER_58_732 ();
 fill_1 FILLER_58_741 ();
 fill_2 FILLER_58_746 ();
 fill_1 FILLER_58_748 ();
 fill_1 FILLER_58_774 ();
 fill_1 FILLER_58_811 ();
 fill_2 FILLER_58_825 ();
 fill_2 FILLER_58_845 ();
 fill_1 FILLER_58_867 ();
 fill_1 FILLER_58_878 ();
 fill_1 FILLER_58_903 ();
 fill_1 FILLER_58_979 ();
 fill_2 FILLER_58_1004 ();
 fill_4 FILLER_58_1013 ();
 fill_1 FILLER_58_1035 ();
 fill_1 FILLER_58_1037 ();
 fill_4 FILLER_59_3 ();
 fill_1 FILLER_59_7 ();
 fill_2 FILLER_59_20 ();
 fill_4 FILLER_59_52 ();
 fill_4 FILLER_59_67 ();
 fill_2 FILLER_59_146 ();
 fill_1 FILLER_59_148 ();
 fill_2 FILLER_59_156 ();
 fill_2 FILLER_59_166 ();
 fill_4 FILLER_59_182 ();
 fill_1 FILLER_59_186 ();
 fill_4 FILLER_59_194 ();
 fill_2 FILLER_59_206 ();
 fill_1 FILLER_59_208 ();
 fill_2 FILLER_59_222 ();
 fill_2 FILLER_59_225 ();
 fill_1 FILLER_59_231 ();
 fill_1 FILLER_59_239 ();
 fill_2 FILLER_59_251 ();
 fill_1 FILLER_59_253 ();
 fill_1 FILLER_59_272 ();
 fill_2 FILLER_59_281 ();
 fill_2 FILLER_59_291 ();
 fill_2 FILLER_59_328 ();
 fill_1 FILLER_59_335 ();
 fill_2 FILLER_59_341 ();
 fill_4 FILLER_59_370 ();
 fill_1 FILLER_59_374 ();
 fill_4 FILLER_59_393 ();
 fill_1 FILLER_59_407 ();
 fill_1 FILLER_59_424 ();
 fill_2 FILLER_59_434 ();
 fill_1 FILLER_59_449 ();
 decap_12 FILLER_59_482 ();
 fill_8 FILLER_59_494 ();
 fill_2 FILLER_59_502 ();
 fill_4 FILLER_59_510 ();
 fill_4 FILLER_59_530 ();
 fill_2 FILLER_59_547 ();
 fill_1 FILLER_59_549 ();
 fill_4 FILLER_59_594 ();
 fill_1 FILLER_59_605 ();
 fill_2 FILLER_59_613 ();
 fill_1 FILLER_59_615 ();
 decap_12 FILLER_59_617 ();
 fill_1 FILLER_59_629 ();
 fill_2 FILLER_59_648 ();
 fill_1 FILLER_59_650 ();
 fill_2 FILLER_59_659 ();
 fill_2 FILLER_59_681 ();
 fill_2 FILLER_59_712 ();
 fill_1 FILLER_59_714 ();
 fill_4 FILLER_59_724 ();
 fill_8 FILLER_59_743 ();
 fill_2 FILLER_59_751 ();
 fill_1 FILLER_59_753 ();
 fill_2 FILLER_59_761 ();
 fill_1 FILLER_59_777 ();
 fill_2 FILLER_59_794 ();
 fill_1 FILLER_59_833 ();
 fill_4 FILLER_59_1004 ();
 fill_2 FILLER_59_1009 ();
 fill_1 FILLER_59_1011 ();
 fill_2 FILLER_60_18 ();
 fill_1 FILLER_60_20 ();
 fill_1 FILLER_60_34 ();
 fill_1 FILLER_60_51 ();
 fill_4 FILLER_60_80 ();
 fill_1 FILLER_60_93 ();
 fill_1 FILLER_60_123 ();
 fill_2 FILLER_60_137 ();
 fill_1 FILLER_60_139 ();
 fill_2 FILLER_60_141 ();
 fill_1 FILLER_60_148 ();
 fill_2 FILLER_60_164 ();
 fill_1 FILLER_60_166 ();
 fill_4 FILLER_60_183 ();
 fill_2 FILLER_60_187 ();
 fill_2 FILLER_60_197 ();
 fill_1 FILLER_60_207 ();
 fill_2 FILLER_60_227 ();
 decap_12 FILLER_60_236 ();
 fill_2 FILLER_60_273 ();
 fill_2 FILLER_60_291 ();
 fill_2 FILLER_60_302 ();
 fill_1 FILLER_60_309 ();
 fill_2 FILLER_60_327 ();
 fill_1 FILLER_60_365 ();
 fill_1 FILLER_60_389 ();
 fill_2 FILLER_60_430 ();
 fill_4 FILLER_60_443 ();
 fill_2 FILLER_60_464 ();
 fill_2 FILLER_60_473 ();
 fill_1 FILLER_60_475 ();
 fill_8 FILLER_60_477 ();
 fill_1 FILLER_60_485 ();
 fill_2 FILLER_60_500 ();
 fill_1 FILLER_60_502 ();
 decap_12 FILLER_60_510 ();
 fill_2 FILLER_60_522 ();
 fill_1 FILLER_60_524 ();
 fill_1 FILLER_60_531 ();
 fill_4 FILLER_60_533 ();
 fill_1 FILLER_60_545 ();
 fill_2 FILLER_60_553 ();
 fill_1 FILLER_60_555 ();
 fill_4 FILLER_60_569 ();
 fill_1 FILLER_60_573 ();
 fill_2 FILLER_60_582 ();
 fill_2 FILLER_60_589 ();
 fill_1 FILLER_60_591 ();
 fill_1 FILLER_60_629 ();
 fill_4 FILLER_60_640 ();
 fill_1 FILLER_60_645 ();
 fill_1 FILLER_60_660 ();
 fill_4 FILLER_60_695 ();
 fill_1 FILLER_60_699 ();
 fill_4 FILLER_60_715 ();
 fill_1 FILLER_60_722 ();
 fill_2 FILLER_60_739 ();
 fill_1 FILLER_60_755 ();
 fill_4 FILLER_60_774 ();
 fill_2 FILLER_60_778 ();
 fill_1 FILLER_60_780 ();
 fill_2 FILLER_60_785 ();
 fill_1 FILLER_60_787 ();
 fill_1 FILLER_60_833 ();
 fill_1 FILLER_60_907 ();
 fill_1 FILLER_60_917 ();
 fill_2 FILLER_60_934 ();
 fill_1 FILLER_60_936 ();
 fill_2 FILLER_60_981 ();
 fill_2 FILLER_60_989 ();
 fill_1 FILLER_60_991 ();
 fill_1 FILLER_60_1037 ();
 fill_1 FILLER_61_3 ();
 fill_1 FILLER_61_23 ();
 fill_1 FILLER_61_34 ();
 fill_2 FILLER_61_45 ();
 fill_1 FILLER_61_47 ();
 fill_4 FILLER_61_70 ();
 fill_4 FILLER_61_108 ();
 fill_4 FILLER_61_113 ();
 fill_4 FILLER_61_122 ();
 decap_12 FILLER_61_130 ();
 fill_2 FILLER_61_142 ();
 fill_1 FILLER_61_148 ();
 fill_4 FILLER_61_163 ();
 fill_1 FILLER_61_167 ();
 fill_2 FILLER_61_169 ();
 fill_2 FILLER_61_175 ();
 fill_8 FILLER_61_207 ();
 fill_1 FILLER_61_215 ();
 fill_2 FILLER_61_221 ();
 fill_1 FILLER_61_223 ();
 fill_4 FILLER_61_225 ();
 fill_4 FILLER_61_236 ();
 fill_4 FILLER_61_268 ();
 fill_2 FILLER_61_281 ();
 fill_2 FILLER_61_291 ();
 fill_1 FILLER_61_293 ();
 fill_2 FILLER_61_341 ();
 fill_1 FILLER_61_343 ();
 fill_2 FILLER_61_358 ();
 fill_1 FILLER_61_360 ();
 fill_1 FILLER_61_364 ();
 fill_4 FILLER_61_376 ();
 fill_2 FILLER_61_380 ();
 fill_1 FILLER_61_382 ();
 fill_1 FILLER_61_387 ();
 fill_8 FILLER_61_410 ();
 fill_2 FILLER_61_445 ();
 fill_1 FILLER_61_447 ();
 decap_12 FILLER_61_488 ();
 fill_4 FILLER_61_500 ();
 fill_4 FILLER_61_505 ();
 fill_2 FILLER_61_509 ();
 decap_12 FILLER_61_518 ();
 decap_12 FILLER_61_530 ();
 decap_12 FILLER_61_542 ();
 fill_4 FILLER_61_554 ();
 fill_2 FILLER_61_558 ();
 fill_2 FILLER_61_567 ();
 fill_1 FILLER_61_569 ();
 fill_8 FILLER_61_586 ();
 fill_1 FILLER_61_594 ();
 fill_1 FILLER_61_602 ();
 fill_4 FILLER_61_612 ();
 fill_1 FILLER_61_617 ();
 fill_8 FILLER_61_645 ();
 fill_1 FILLER_61_653 ();
 fill_4 FILLER_61_691 ();
 fill_2 FILLER_61_695 ();
 fill_4 FILLER_61_708 ();
 fill_2 FILLER_61_719 ();
 decap_12 FILLER_61_729 ();
 decap_12 FILLER_61_741 ();
 decap_12 FILLER_61_753 ();
 fill_4 FILLER_61_765 ();
 fill_8 FILLER_61_776 ();
 fill_2 FILLER_61_794 ();
 fill_1 FILLER_61_796 ();
 fill_4 FILLER_61_800 ();
 fill_2 FILLER_61_804 ();
 fill_2 FILLER_61_809 ();
 fill_2 FILLER_61_817 ();
 fill_2 FILLER_61_838 ();
 fill_1 FILLER_61_850 ();
 fill_1 FILLER_61_872 ();
 fill_1 FILLER_61_917 ();
 fill_1 FILLER_61_941 ();
 fill_1 FILLER_61_951 ();
 fill_1 FILLER_61_965 ();
 fill_1 FILLER_61_1004 ();
 fill_4 FILLER_62_23 ();
 fill_1 FILLER_62_27 ();
 fill_1 FILLER_62_29 ();
 fill_1 FILLER_62_41 ();
 fill_2 FILLER_62_77 ();
 fill_1 FILLER_62_93 ();
 fill_1 FILLER_62_101 ();
 fill_1 FILLER_62_110 ();
 fill_2 FILLER_62_130 ();
 fill_2 FILLER_62_141 ();
 fill_1 FILLER_62_143 ();
 fill_1 FILLER_62_148 ();
 decap_12 FILLER_62_155 ();
 fill_2 FILLER_62_167 ();
 fill_2 FILLER_62_176 ();
 fill_1 FILLER_62_178 ();
 fill_1 FILLER_62_188 ();
 fill_1 FILLER_62_197 ();
 fill_1 FILLER_62_210 ();
 fill_8 FILLER_62_225 ();
 fill_4 FILLER_62_240 ();
 fill_1 FILLER_62_244 ();
 fill_2 FILLER_62_253 ();
 fill_4 FILLER_62_270 ();
 fill_1 FILLER_62_274 ();
 fill_1 FILLER_62_309 ();
 fill_2 FILLER_62_322 ();
 fill_4 FILLER_62_331 ();
 fill_1 FILLER_62_335 ();
 fill_2 FILLER_62_362 ();
 fill_2 FILLER_62_365 ();
 fill_2 FILLER_62_379 ();
 fill_2 FILLER_62_411 ();
 fill_8 FILLER_62_466 ();
 fill_2 FILLER_62_474 ();
 fill_4 FILLER_62_477 ();
 fill_1 FILLER_62_481 ();
 fill_4 FILLER_62_489 ();
 fill_1 FILLER_62_493 ();
 fill_8 FILLER_62_504 ();
 decap_12 FILLER_62_519 ();
 fill_1 FILLER_62_531 ();
 decap_12 FILLER_62_533 ();
 fill_8 FILLER_62_545 ();
 fill_8 FILLER_62_568 ();
 fill_1 FILLER_62_576 ();
 fill_2 FILLER_62_586 ();
 fill_2 FILLER_62_599 ();
 fill_1 FILLER_62_601 ();
 decap_12 FILLER_62_619 ();
 decap_12 FILLER_62_631 ();
 fill_1 FILLER_62_643 ();
 fill_2 FILLER_62_662 ();
 fill_1 FILLER_62_664 ();
 fill_2 FILLER_62_697 ();
 fill_1 FILLER_62_699 ();
 fill_2 FILLER_62_715 ();
 fill_1 FILLER_62_717 ();
 fill_2 FILLER_62_764 ();
 decap_12 FILLER_62_773 ();
 fill_2 FILLER_62_800 ();
 fill_1 FILLER_62_802 ();
 fill_2 FILLER_62_819 ();
 fill_1 FILLER_62_844 ();
 fill_1 FILLER_62_902 ();
 fill_2 FILLER_62_921 ();
 fill_1 FILLER_62_923 ();
 fill_2 FILLER_62_925 ();
 fill_2 FILLER_62_968 ();
 fill_1 FILLER_62_970 ();
 fill_2 FILLER_62_1010 ();
 fill_1 FILLER_62_1012 ();
 fill_1 FILLER_62_1022 ();
 fill_1 FILLER_62_1035 ();
 fill_1 FILLER_62_1037 ();
 fill_4 FILLER_63_30 ();
 fill_2 FILLER_63_34 ();
 fill_2 FILLER_63_76 ();
 fill_1 FILLER_63_78 ();
 fill_1 FILLER_63_90 ();
 fill_2 FILLER_63_110 ();
 fill_4 FILLER_63_120 ();
 fill_8 FILLER_63_140 ();
 fill_4 FILLER_63_156 ();
 fill_1 FILLER_63_160 ();
 fill_2 FILLER_63_180 ();
 fill_1 FILLER_63_182 ();
 fill_8 FILLER_63_200 ();
 fill_2 FILLER_63_208 ();
 fill_1 FILLER_63_210 ();
 fill_8 FILLER_63_214 ();
 fill_2 FILLER_63_222 ();
 decap_12 FILLER_63_232 ();
 decap_12 FILLER_63_244 ();
 fill_4 FILLER_63_256 ();
 fill_2 FILLER_63_260 ();
 fill_2 FILLER_63_323 ();
 fill_1 FILLER_63_325 ();
 fill_1 FILLER_63_342 ();
 fill_1 FILLER_63_369 ();
 decap_12 FILLER_63_374 ();
 fill_1 FILLER_63_393 ();
 fill_2 FILLER_63_446 ();
 fill_2 FILLER_63_474 ();
 fill_1 FILLER_63_476 ();
 fill_4 FILLER_63_483 ();
 fill_2 FILLER_63_487 ();
 fill_4 FILLER_63_497 ();
 fill_2 FILLER_63_501 ();
 fill_1 FILLER_63_503 ();
 fill_4 FILLER_63_549 ();
 fill_2 FILLER_63_553 ();
 fill_2 FILLER_63_558 ();
 fill_2 FILLER_63_566 ();
 fill_8 FILLER_63_582 ();
 decap_12 FILLER_63_593 ();
 fill_8 FILLER_63_605 ();
 fill_2 FILLER_63_613 ();
 fill_1 FILLER_63_615 ();
 fill_2 FILLER_63_634 ();
 fill_1 FILLER_63_653 ();
 fill_2 FILLER_63_670 ();
 fill_8 FILLER_63_686 ();
 fill_2 FILLER_63_701 ();
 decap_12 FILLER_63_711 ();
 fill_4 FILLER_63_723 ();
 fill_1 FILLER_63_727 ();
 fill_8 FILLER_63_729 ();
 fill_2 FILLER_63_737 ();
 fill_2 FILLER_63_782 ();
 fill_2 FILLER_63_825 ();
 fill_1 FILLER_63_827 ();
 fill_2 FILLER_63_837 ();
 fill_1 FILLER_63_839 ();
 fill_2 FILLER_63_841 ();
 fill_1 FILLER_63_892 ();
 fill_4 FILLER_63_906 ();
 fill_2 FILLER_63_910 ();
 fill_1 FILLER_63_912 ();
 fill_4 FILLER_63_936 ();
 fill_1 FILLER_63_940 ();
 fill_1 FILLER_63_951 ();
 fill_8 FILLER_63_980 ();
 fill_2 FILLER_63_988 ();
 fill_2 FILLER_63_1005 ();
 fill_1 FILLER_63_1007 ();
 fill_2 FILLER_64_3 ();
 fill_1 FILLER_64_5 ();
 fill_2 FILLER_64_13 ();
 fill_8 FILLER_64_20 ();
 fill_1 FILLER_64_29 ();
 fill_8 FILLER_64_37 ();
 fill_4 FILLER_64_60 ();
 fill_1 FILLER_64_83 ();
 fill_4 FILLER_64_85 ();
 fill_4 FILLER_64_145 ();
 fill_2 FILLER_64_154 ();
 fill_1 FILLER_64_208 ();
 fill_4 FILLER_64_221 ();
 fill_4 FILLER_64_233 ();
 fill_2 FILLER_64_237 ();
 fill_1 FILLER_64_239 ();
 fill_4 FILLER_64_248 ();
 fill_8 FILLER_64_253 ();
 fill_1 FILLER_64_261 ();
 fill_4 FILLER_64_284 ();
 fill_2 FILLER_64_288 ();
 fill_2 FILLER_64_306 ();
 fill_1 FILLER_64_340 ();
 fill_4 FILLER_64_358 ();
 fill_2 FILLER_64_362 ();
 fill_8 FILLER_64_365 ();
 fill_1 FILLER_64_373 ();
 fill_2 FILLER_64_456 ();
 fill_1 FILLER_64_458 ();
 fill_4 FILLER_64_462 ();
 fill_2 FILLER_64_466 ();
 fill_1 FILLER_64_468 ();
 decap_12 FILLER_64_502 ();
 fill_4 FILLER_64_514 ();
 fill_1 FILLER_64_518 ();
 fill_1 FILLER_64_531 ();
 decap_12 FILLER_64_533 ();
 decap_12 FILLER_64_545 ();
 fill_1 FILLER_64_557 ();
 fill_4 FILLER_64_567 ();
 fill_2 FILLER_64_571 ();
 fill_1 FILLER_64_573 ();
 fill_2 FILLER_64_585 ();
 fill_1 FILLER_64_587 ();
 fill_2 FILLER_64_596 ();
 fill_1 FILLER_64_622 ();
 fill_1 FILLER_64_627 ();
 fill_1 FILLER_64_643 ();
 fill_4 FILLER_64_645 ();
 fill_2 FILLER_64_649 ();
 decap_12 FILLER_64_663 ();
 fill_4 FILLER_64_675 ();
 fill_1 FILLER_64_679 ();
 fill_4 FILLER_64_687 ();
 fill_2 FILLER_64_691 ();
 fill_1 FILLER_64_693 ();
 fill_1 FILLER_64_704 ();
 fill_8 FILLER_64_715 ();
 fill_1 FILLER_64_739 ();
 fill_1 FILLER_64_743 ();
 fill_8 FILLER_64_747 ();
 fill_1 FILLER_64_755 ();
 decap_12 FILLER_64_764 ();
 fill_1 FILLER_64_776 ();
 fill_4 FILLER_64_784 ();
 fill_2 FILLER_64_788 ();
 fill_1 FILLER_64_790 ();
 fill_2 FILLER_64_804 ();
 fill_2 FILLER_64_826 ();
 fill_1 FILLER_64_854 ();
 fill_4 FILLER_64_864 ();
 fill_4 FILLER_64_869 ();
 fill_2 FILLER_64_882 ();
 fill_2 FILLER_64_907 ();
 fill_1 FILLER_64_909 ();
 fill_4 FILLER_64_919 ();
 fill_1 FILLER_64_923 ();
 fill_2 FILLER_64_940 ();
 fill_1 FILLER_64_942 ();
 fill_2 FILLER_64_949 ();
 fill_1 FILLER_64_951 ();
 fill_2 FILLER_64_956 ();
 fill_2 FILLER_64_978 ();
 fill_4 FILLER_64_981 ();
 fill_2 FILLER_64_1009 ();
 fill_2 FILLER_64_1017 ();
 fill_1 FILLER_64_1019 ();
 fill_1 FILLER_64_1032 ();
 fill_1 FILLER_64_1037 ();
 fill_4 FILLER_65_3 ();
 fill_1 FILLER_65_7 ();
 fill_1 FILLER_65_20 ();
 fill_2 FILLER_65_44 ();
 fill_1 FILLER_65_46 ();
 fill_2 FILLER_65_57 ();
 fill_2 FILLER_65_97 ();
 fill_1 FILLER_65_99 ();
 fill_2 FILLER_65_116 ();
 fill_1 FILLER_65_118 ();
 decap_12 FILLER_65_123 ();
 fill_8 FILLER_65_135 ();
 fill_2 FILLER_65_185 ();
 fill_2 FILLER_65_204 ();
 fill_1 FILLER_65_206 ();
 fill_4 FILLER_65_220 ();
 fill_1 FILLER_65_232 ();
 fill_2 FILLER_65_278 ();
 fill_4 FILLER_65_281 ();
 fill_2 FILLER_65_285 ();
 fill_2 FILLER_65_304 ();
 fill_2 FILLER_65_328 ();
 fill_4 FILLER_65_343 ();
 fill_2 FILLER_65_347 ();
 fill_1 FILLER_65_375 ();
 fill_4 FILLER_65_409 ();
 fill_1 FILLER_65_429 ();
 fill_2 FILLER_65_446 ();
 fill_2 FILLER_65_449 ();
 fill_1 FILLER_65_460 ();
 fill_2 FILLER_65_466 ();
 fill_1 FILLER_65_468 ();
 fill_4 FILLER_65_484 ();
 fill_1 FILLER_65_503 ();
 fill_2 FILLER_65_520 ();
 fill_2 FILLER_65_531 ();
 fill_1 FILLER_65_533 ();
 fill_1 FILLER_65_559 ();
 fill_1 FILLER_65_592 ();
 fill_4 FILLER_65_609 ();
 fill_2 FILLER_65_613 ();
 fill_1 FILLER_65_615 ();
 fill_2 FILLER_65_617 ();
 fill_1 FILLER_65_619 ();
 decap_12 FILLER_65_631 ();
 fill_2 FILLER_65_643 ();
 fill_1 FILLER_65_645 ();
 fill_2 FILLER_65_670 ();
 fill_8 FILLER_65_680 ();
 fill_1 FILLER_65_704 ();
 fill_4 FILLER_65_722 ();
 fill_2 FILLER_65_726 ();
 fill_8 FILLER_65_729 ();
 fill_2 FILLER_65_737 ();
 fill_1 FILLER_65_747 ();
 fill_4 FILLER_65_755 ();
 fill_2 FILLER_65_759 ();
 fill_4 FILLER_65_778 ();
 fill_2 FILLER_65_782 ();
 fill_2 FILLER_65_805 ();
 fill_1 FILLER_65_807 ();
 fill_1 FILLER_65_853 ();
 fill_4 FILLER_65_860 ();
 fill_1 FILLER_65_887 ();
 fill_2 FILLER_65_894 ();
 fill_4 FILLER_65_915 ();
 fill_2 FILLER_65_919 ();
 fill_1 FILLER_65_921 ();
 fill_1 FILLER_65_988 ();
 fill_1 FILLER_65_1004 ();
 fill_1 FILLER_65_1009 ();
 fill_2 FILLER_65_1036 ();
 fill_1 FILLER_66_27 ();
 fill_4 FILLER_66_29 ();
 fill_8 FILLER_66_39 ();
 fill_2 FILLER_66_55 ();
 fill_4 FILLER_66_85 ();
 fill_2 FILLER_66_89 ();
 fill_1 FILLER_66_91 ();
 fill_1 FILLER_66_108 ();
 fill_1 FILLER_66_122 ();
 fill_2 FILLER_66_131 ();
 fill_2 FILLER_66_138 ();
 fill_2 FILLER_66_150 ();
 fill_2 FILLER_66_197 ();
 decap_12 FILLER_66_225 ();
 decap_12 FILLER_66_237 ();
 fill_2 FILLER_66_249 ();
 fill_1 FILLER_66_251 ();
 decap_12 FILLER_66_253 ();
 fill_2 FILLER_66_265 ();
 fill_1 FILLER_66_267 ();
 fill_4 FILLER_66_292 ();
 fill_1 FILLER_66_296 ();
 fill_2 FILLER_66_318 ();
 fill_1 FILLER_66_356 ();
 fill_1 FILLER_66_363 ();
 fill_8 FILLER_66_365 ();
 fill_1 FILLER_66_373 ();
 fill_8 FILLER_66_389 ();
 fill_2 FILLER_66_397 ();
 fill_1 FILLER_66_399 ();
 fill_4 FILLER_66_407 ();
 fill_2 FILLER_66_418 ();
 fill_1 FILLER_66_443 ();
 fill_4 FILLER_66_471 ();
 fill_1 FILLER_66_475 ();
 fill_2 FILLER_66_477 ();
 fill_4 FILLER_66_496 ();
 fill_1 FILLER_66_516 ();
 fill_2 FILLER_66_523 ();
 fill_2 FILLER_66_530 ();
 fill_4 FILLER_66_533 ();
 fill_1 FILLER_66_537 ();
 fill_4 FILLER_66_544 ();
 fill_1 FILLER_66_555 ();
 fill_8 FILLER_66_565 ();
 fill_1 FILLER_66_573 ();
 fill_4 FILLER_66_581 ();
 fill_2 FILLER_66_585 ();
 fill_1 FILLER_66_587 ();
 fill_2 FILLER_66_598 ();
 fill_1 FILLER_66_600 ();
 fill_4 FILLER_66_633 ();
 fill_1 FILLER_66_645 ();
 fill_4 FILLER_66_653 ();
 fill_2 FILLER_66_657 ();
 fill_2 FILLER_66_666 ();
 fill_1 FILLER_66_668 ();
 fill_1 FILLER_66_699 ();
 fill_4 FILLER_66_708 ();
 fill_2 FILLER_66_712 ();
 fill_1 FILLER_66_736 ();
 fill_2 FILLER_66_754 ();
 fill_4 FILLER_66_764 ();
 fill_2 FILLER_66_768 ();
 fill_1 FILLER_66_770 ();
 fill_8 FILLER_66_781 ();
 fill_1 FILLER_66_789 ();
 fill_1 FILLER_66_811 ();
 fill_2 FILLER_66_816 ();
 fill_2 FILLER_66_836 ();
 fill_2 FILLER_66_847 ();
 fill_2 FILLER_66_869 ();
 fill_1 FILLER_66_871 ();
 fill_2 FILLER_66_888 ();
 fill_1 FILLER_66_923 ();
 fill_1 FILLER_66_990 ();
 fill_4 FILLER_66_1000 ();
 fill_2 FILLER_66_1025 ();
 fill_1 FILLER_66_1027 ();
 fill_4 FILLER_66_1031 ();
 fill_1 FILLER_66_1035 ();
 fill_1 FILLER_66_1037 ();
 fill_4 FILLER_67_3 ();
 fill_2 FILLER_67_7 ();
 fill_1 FILLER_67_24 ();
 fill_1 FILLER_67_42 ();
 fill_1 FILLER_67_55 ();
 fill_1 FILLER_67_60 ();
 fill_4 FILLER_67_69 ();
 fill_1 FILLER_67_73 ();
 fill_1 FILLER_67_94 ();
 fill_2 FILLER_67_113 ();
 fill_2 FILLER_67_135 ();
 fill_4 FILLER_67_148 ();
 fill_1 FILLER_67_158 ();
 fill_1 FILLER_67_183 ();
 fill_2 FILLER_67_221 ();
 fill_1 FILLER_67_223 ();
 fill_1 FILLER_67_244 ();
 fill_1 FILLER_67_252 ();
 fill_4 FILLER_67_265 ();
 fill_4 FILLER_67_276 ();
 fill_1 FILLER_67_296 ();
 fill_8 FILLER_67_301 ();
 fill_2 FILLER_67_313 ();
 fill_1 FILLER_67_337 ();
 fill_2 FILLER_67_349 ();
 fill_2 FILLER_67_390 ();
 fill_4 FILLER_67_397 ();
 fill_1 FILLER_67_418 ();
 fill_2 FILLER_67_445 ();
 fill_1 FILLER_67_447 ();
 fill_1 FILLER_67_452 ();
 fill_4 FILLER_67_461 ();
 fill_1 FILLER_67_480 ();
 fill_2 FILLER_67_488 ();
 fill_1 FILLER_67_490 ();
 fill_4 FILLER_67_499 ();
 fill_1 FILLER_67_503 ();
 fill_2 FILLER_67_521 ();
 fill_1 FILLER_67_523 ();
 fill_2 FILLER_67_530 ();
 fill_1 FILLER_67_532 ();
 fill_2 FILLER_67_541 ();
 fill_1 FILLER_67_543 ();
 fill_2 FILLER_67_550 ();
 fill_1 FILLER_67_565 ();
 fill_2 FILLER_67_596 ();
 fill_1 FILLER_67_598 ();
 fill_4 FILLER_67_609 ();
 fill_2 FILLER_67_613 ();
 fill_1 FILLER_67_615 ();
 fill_4 FILLER_67_626 ();
 fill_2 FILLER_67_630 ();
 fill_2 FILLER_67_652 ();
 fill_2 FILLER_67_670 ();
 fill_2 FILLER_67_680 ();
 fill_1 FILLER_67_682 ();
 fill_2 FILLER_67_691 ();
 fill_1 FILLER_67_693 ();
 decap_12 FILLER_67_701 ();
 fill_2 FILLER_67_713 ();
 fill_2 FILLER_67_722 ();
 fill_1 FILLER_67_724 ();
 fill_2 FILLER_67_737 ();
 fill_4 FILLER_67_748 ();
 fill_4 FILLER_67_755 ();
 fill_1 FILLER_67_769 ();
 fill_2 FILLER_67_782 ();
 fill_1 FILLER_67_830 ();
 fill_1 FILLER_67_897 ();
 fill_2 FILLER_67_907 ();
 fill_1 FILLER_67_909 ();
 fill_1 FILLER_67_922 ();
 fill_2 FILLER_67_950 ();
 fill_2 FILLER_67_985 ();
 fill_1 FILLER_67_1007 ();
 fill_2 FILLER_67_1036 ();
 fill_1 FILLER_68_27 ();
 fill_1 FILLER_68_29 ();
 fill_1 FILLER_68_50 ();
 fill_1 FILLER_68_78 ();
 fill_2 FILLER_68_85 ();
 fill_1 FILLER_68_98 ();
 fill_4 FILLER_68_106 ();
 fill_8 FILLER_68_130 ();
 fill_2 FILLER_68_138 ();
 fill_2 FILLER_68_170 ();
 fill_1 FILLER_68_195 ();
 decap_12 FILLER_68_217 ();
 fill_2 FILLER_68_229 ();
 fill_4 FILLER_68_238 ();
 fill_1 FILLER_68_242 ();
 fill_2 FILLER_68_250 ();
 fill_4 FILLER_68_260 ();
 fill_1 FILLER_68_264 ();
 fill_1 FILLER_68_282 ();
 fill_1 FILLER_68_302 ();
 fill_2 FILLER_68_318 ();
 fill_1 FILLER_68_356 ();
 fill_1 FILLER_68_363 ();
 fill_1 FILLER_68_365 ();
 fill_1 FILLER_68_374 ();
 fill_4 FILLER_68_408 ();
 fill_1 FILLER_68_412 ();
 fill_2 FILLER_68_421 ();
 fill_1 FILLER_68_432 ();
 fill_4 FILLER_68_441 ();
 fill_1 FILLER_68_484 ();
 fill_4 FILLER_68_494 ();
 fill_1 FILLER_68_498 ();
 fill_2 FILLER_68_508 ();
 fill_4 FILLER_68_517 ();
 fill_2 FILLER_68_529 ();
 fill_1 FILLER_68_531 ();
 fill_2 FILLER_68_545 ();
 fill_1 FILLER_68_547 ();
 fill_4 FILLER_68_565 ();
 fill_1 FILLER_68_569 ();
 decap_12 FILLER_68_576 ();
 fill_4 FILLER_68_609 ();
 fill_8 FILLER_68_630 ();
 fill_2 FILLER_68_638 ();
 fill_1 FILLER_68_640 ();
 fill_2 FILLER_68_645 ();
 fill_2 FILLER_68_659 ();
 fill_1 FILLER_68_661 ();
 fill_8 FILLER_68_669 ();
 decap_12 FILLER_68_684 ();
 fill_4 FILLER_68_696 ();
 fill_4 FILLER_68_701 ();
 fill_1 FILLER_68_712 ();
 fill_2 FILLER_68_754 ();
 fill_2 FILLER_68_769 ();
 fill_4 FILLER_68_778 ();
 fill_2 FILLER_68_782 ();
 fill_1 FILLER_68_784 ();
 fill_1 FILLER_68_811 ();
 fill_4 FILLER_68_813 ();
 fill_2 FILLER_68_817 ();
 fill_1 FILLER_68_819 ();
 fill_4 FILLER_68_829 ();
 fill_2 FILLER_68_845 ();
 fill_1 FILLER_68_847 ();
 fill_4 FILLER_68_863 ();
 fill_1 FILLER_68_867 ();
 fill_2 FILLER_68_872 ();
 fill_1 FILLER_68_874 ();
 fill_2 FILLER_68_948 ();
 fill_1 FILLER_68_981 ();
 fill_2 FILLER_68_997 ();
 fill_4 FILLER_68_1008 ();
 fill_1 FILLER_68_1012 ();
 fill_1 FILLER_68_1037 ();
 fill_8 FILLER_69_3 ();
 fill_2 FILLER_69_20 ();
 fill_2 FILLER_69_25 ();
 fill_2 FILLER_69_38 ();
 fill_8 FILLER_69_45 ();
 fill_4 FILLER_69_62 ();
 fill_2 FILLER_69_66 ();
 fill_1 FILLER_69_68 ();
 fill_2 FILLER_69_77 ();
 fill_1 FILLER_69_113 ();
 fill_2 FILLER_69_140 ();
 fill_2 FILLER_69_156 ();
 fill_1 FILLER_69_167 ();
 fill_1 FILLER_69_178 ();
 fill_1 FILLER_69_214 ();
 fill_2 FILLER_69_222 ();
 decap_12 FILLER_69_225 ();
 fill_1 FILLER_69_237 ();
 fill_2 FILLER_69_243 ();
 decap_12 FILLER_69_252 ();
 fill_4 FILLER_69_264 ();
 fill_4 FILLER_69_275 ();
 fill_1 FILLER_69_279 ();
 fill_1 FILLER_69_285 ();
 fill_1 FILLER_69_300 ();
 fill_2 FILLER_69_334 ();
 fill_2 FILLER_69_343 ();
 fill_1 FILLER_69_345 ();
 fill_4 FILLER_69_425 ();
 fill_2 FILLER_69_437 ();
 fill_2 FILLER_69_446 ();
 fill_4 FILLER_69_457 ();
 decap_12 FILLER_69_492 ();
 fill_4 FILLER_69_505 ();
 fill_2 FILLER_69_517 ();
 fill_2 FILLER_69_527 ();
 fill_1 FILLER_69_529 ();
 fill_2 FILLER_69_538 ();
 fill_4 FILLER_69_556 ();
 fill_2 FILLER_69_561 ();
 fill_1 FILLER_69_563 ();
 fill_2 FILLER_69_571 ();
 fill_1 FILLER_69_573 ();
 fill_4 FILLER_69_588 ();
 fill_2 FILLER_69_592 ();
 fill_1 FILLER_69_594 ();
 fill_4 FILLER_69_602 ();
 fill_2 FILLER_69_606 ();
 fill_1 FILLER_69_615 ();
 fill_4 FILLER_69_617 ();
 fill_2 FILLER_69_631 ();
 fill_1 FILLER_69_633 ();
 fill_2 FILLER_69_641 ();
 fill_2 FILLER_69_650 ();
 fill_1 FILLER_69_652 ();
 fill_8 FILLER_69_662 ();
 fill_2 FILLER_69_670 ();
 fill_1 FILLER_69_680 ();
 fill_1 FILLER_69_702 ();
 fill_2 FILLER_69_710 ();
 fill_4 FILLER_69_718 ();
 fill_2 FILLER_69_722 ();
 fill_1 FILLER_69_724 ();
 fill_2 FILLER_69_738 ();
 fill_4 FILLER_69_747 ();
 fill_2 FILLER_69_751 ();
 fill_1 FILLER_69_765 ();
 fill_8 FILLER_69_773 ();
 fill_2 FILLER_69_781 ();
 fill_1 FILLER_69_783 ();
 fill_8 FILLER_69_801 ();
 fill_2 FILLER_69_809 ();
 fill_2 FILLER_69_838 ();
 fill_1 FILLER_69_861 ();
 fill_1 FILLER_69_895 ();
 fill_2 FILLER_69_903 ();
 fill_2 FILLER_69_929 ();
 fill_1 FILLER_69_931 ();
 fill_2 FILLER_69_962 ();
 fill_1 FILLER_69_1007 ();
 fill_4 FILLER_69_1009 ();
 fill_1 FILLER_69_1013 ();
 fill_1 FILLER_69_1020 ();
 fill_8 FILLER_69_1030 ();
 fill_1 FILLER_70_20 ();
 fill_1 FILLER_70_45 ();
 fill_2 FILLER_70_81 ();
 fill_1 FILLER_70_83 ();
 fill_2 FILLER_70_85 ();
 fill_1 FILLER_70_87 ();
 fill_4 FILLER_70_95 ();
 fill_2 FILLER_70_112 ();
 fill_1 FILLER_70_114 ();
 fill_2 FILLER_70_138 ();
 fill_1 FILLER_70_165 ();
 decap_12 FILLER_70_206 ();
 fill_8 FILLER_70_218 ();
 fill_8 FILLER_70_236 ();
 fill_1 FILLER_70_244 ();
 fill_4 FILLER_70_274 ();
 fill_8 FILLER_70_298 ();
 fill_2 FILLER_70_306 ();
 fill_2 FILLER_70_314 ();
 fill_2 FILLER_70_322 ();
 fill_2 FILLER_70_347 ();
 fill_2 FILLER_70_362 ();
 fill_8 FILLER_70_368 ();
 fill_2 FILLER_70_376 ();
 fill_4 FILLER_70_386 ();
 fill_2 FILLER_70_390 ();
 fill_2 FILLER_70_412 ();
 fill_1 FILLER_70_414 ();
 fill_2 FILLER_70_421 ();
 fill_1 FILLER_70_423 ();
 fill_4 FILLER_70_458 ();
 fill_2 FILLER_70_474 ();
 fill_4 FILLER_70_477 ();
 fill_4 FILLER_70_505 ();
 fill_4 FILLER_70_521 ();
 fill_2 FILLER_70_525 ();
 fill_1 FILLER_70_531 ();
 decap_12 FILLER_70_533 ();
 fill_4 FILLER_70_545 ();
 fill_8 FILLER_70_561 ();
 fill_2 FILLER_70_569 ();
 fill_8 FILLER_70_577 ();
 fill_2 FILLER_70_585 ();
 fill_1 FILLER_70_587 ();
 decap_12 FILLER_70_596 ();
 decap_12 FILLER_70_608 ();
 fill_2 FILLER_70_626 ();
 fill_1 FILLER_70_628 ();
 fill_8 FILLER_70_636 ();
 fill_4 FILLER_70_645 ();
 fill_1 FILLER_70_649 ();
 fill_2 FILLER_70_667 ();
 fill_1 FILLER_70_669 ();
 fill_8 FILLER_70_678 ();
 fill_2 FILLER_70_686 ();
 fill_4 FILLER_70_695 ();
 fill_1 FILLER_70_699 ();
 fill_4 FILLER_70_701 ();
 fill_2 FILLER_70_705 ();
 fill_1 FILLER_70_707 ();
 fill_4 FILLER_70_715 ();
 fill_2 FILLER_70_726 ();
 fill_1 FILLER_70_731 ();
 fill_4 FILLER_70_757 ();
 fill_1 FILLER_70_761 ();
 fill_8 FILLER_70_769 ();
 fill_1 FILLER_70_777 ();
 fill_4 FILLER_70_807 ();
 fill_1 FILLER_70_811 ();
 fill_2 FILLER_70_822 ();
 fill_2 FILLER_70_856 ();
 fill_1 FILLER_70_858 ();
 fill_1 FILLER_70_878 ();
 fill_2 FILLER_70_894 ();
 fill_4 FILLER_70_905 ();
 fill_1 FILLER_70_909 ();
 fill_4 FILLER_70_913 ();
 fill_1 FILLER_70_917 ();
 fill_4 FILLER_70_934 ();
 fill_1 FILLER_70_938 ();
 fill_1 FILLER_70_971 ();
 fill_2 FILLER_70_978 ();
 fill_4 FILLER_70_981 ();
 fill_1 FILLER_70_985 ();
 fill_1 FILLER_70_1015 ();
 fill_1 FILLER_70_1037 ();
 fill_4 FILLER_71_3 ();
 fill_2 FILLER_71_7 ();
 fill_1 FILLER_71_23 ();
 fill_2 FILLER_71_37 ();
 fill_1 FILLER_71_55 ();
 fill_4 FILLER_71_62 ();
 fill_2 FILLER_71_66 ();
 fill_2 FILLER_71_86 ();
 fill_1 FILLER_71_88 ();
 fill_1 FILLER_71_113 ();
 fill_2 FILLER_71_131 ();
 fill_2 FILLER_71_203 ();
 fill_4 FILLER_71_217 ();
 fill_2 FILLER_71_221 ();
 fill_1 FILLER_71_223 ();
 fill_1 FILLER_71_232 ();
 decap_12 FILLER_71_248 ();
 fill_1 FILLER_71_260 ();
 fill_4 FILLER_71_265 ();
 fill_4 FILLER_71_281 ();
 fill_2 FILLER_71_285 ();
 fill_2 FILLER_71_361 ();
 fill_1 FILLER_71_363 ();
 fill_2 FILLER_71_367 ();
 fill_2 FILLER_71_389 ();
 fill_1 FILLER_71_391 ();
 fill_1 FILLER_71_407 ();
 fill_2 FILLER_71_433 ();
 fill_1 FILLER_71_435 ();
 fill_2 FILLER_71_445 ();
 fill_1 FILLER_71_447 ();
 fill_1 FILLER_71_463 ();
 fill_2 FILLER_71_472 ();
 fill_1 FILLER_71_474 ();
 fill_4 FILLER_71_492 ();
 fill_1 FILLER_71_503 ();
 fill_1 FILLER_71_516 ();
 fill_2 FILLER_71_541 ();
 fill_1 FILLER_71_559 ();
 fill_2 FILLER_71_610 ();
 fill_2 FILLER_71_631 ();
 fill_1 FILLER_71_633 ();
 fill_4 FILLER_71_647 ();
 fill_2 FILLER_71_651 ();
 fill_8 FILLER_71_656 ();
 fill_2 FILLER_71_664 ();
 fill_1 FILLER_71_666 ();
 fill_4 FILLER_71_697 ();
 fill_1 FILLER_71_701 ();
 fill_2 FILLER_71_736 ();
 fill_2 FILLER_71_745 ();
 fill_2 FILLER_71_761 ();
 fill_1 FILLER_71_763 ();
 fill_2 FILLER_71_781 ();
 fill_1 FILLER_71_783 ();
 fill_1 FILLER_71_839 ();
 decap_12 FILLER_71_859 ();
 fill_2 FILLER_71_894 ();
 fill_2 FILLER_71_917 ();
 fill_1 FILLER_71_942 ();
 fill_2 FILLER_71_968 ();
 fill_1 FILLER_71_990 ();
 fill_4 FILLER_71_1000 ();
 fill_1 FILLER_71_1004 ();
 fill_8 FILLER_71_1030 ();
 decap_12 FILLER_72_3 ();
 fill_2 FILLER_72_15 ();
 fill_1 FILLER_72_20 ();
 fill_2 FILLER_72_76 ();
 fill_4 FILLER_72_85 ();
 fill_2 FILLER_72_106 ();
 fill_1 FILLER_72_108 ();
 fill_1 FILLER_72_115 ();
 fill_2 FILLER_72_128 ();
 fill_1 FILLER_72_139 ();
 fill_2 FILLER_72_141 ();
 fill_2 FILLER_72_169 ();
 fill_1 FILLER_72_195 ();
 fill_1 FILLER_72_210 ();
 fill_4 FILLER_72_220 ();
 fill_1 FILLER_72_233 ();
 fill_4 FILLER_72_253 ();
 fill_2 FILLER_72_273 ();
 fill_1 FILLER_72_289 ();
 fill_4 FILLER_72_303 ();
 fill_1 FILLER_72_307 ();
 fill_2 FILLER_72_309 ();
 fill_2 FILLER_72_319 ();
 fill_2 FILLER_72_345 ();
 fill_2 FILLER_72_381 ();
 fill_2 FILLER_72_417 ();
 fill_1 FILLER_72_419 ();
 fill_1 FILLER_72_421 ();
 fill_8 FILLER_72_438 ();
 fill_2 FILLER_72_454 ();
 fill_2 FILLER_72_488 ();
 fill_1 FILLER_72_490 ();
 fill_8 FILLER_72_521 ();
 fill_2 FILLER_72_529 ();
 fill_1 FILLER_72_531 ();
 decap_12 FILLER_72_542 ();
 decap_12 FILLER_72_554 ();
 fill_4 FILLER_72_566 ();
 fill_1 FILLER_72_570 ();
 fill_8 FILLER_72_578 ();
 fill_2 FILLER_72_586 ();
 fill_8 FILLER_72_589 ();
 fill_2 FILLER_72_597 ();
 fill_1 FILLER_72_599 ();
 fill_8 FILLER_72_607 ();
 fill_2 FILLER_72_615 ();
 fill_1 FILLER_72_617 ();
 fill_8 FILLER_72_627 ();
 fill_1 FILLER_72_635 ();
 fill_1 FILLER_72_643 ();
 fill_4 FILLER_72_645 ();
 fill_1 FILLER_72_649 ();
 fill_1 FILLER_72_670 ();
 fill_8 FILLER_72_674 ();
 fill_1 FILLER_72_682 ();
 fill_4 FILLER_72_687 ();
 fill_2 FILLER_72_691 ();
 fill_1 FILLER_72_693 ();
 fill_2 FILLER_72_715 ();
 fill_2 FILLER_72_740 ();
 fill_4 FILLER_72_757 ();
 fill_2 FILLER_72_761 ();
 fill_1 FILLER_72_763 ();
 fill_4 FILLER_72_774 ();
 fill_2 FILLER_72_778 ();
 fill_4 FILLER_72_798 ();
 fill_4 FILLER_72_808 ();
 fill_1 FILLER_72_813 ();
 fill_2 FILLER_72_863 ();
 fill_2 FILLER_72_878 ();
 fill_1 FILLER_72_880 ();
 fill_2 FILLER_72_890 ();
 fill_1 FILLER_72_892 ();
 fill_2 FILLER_72_908 ();
 fill_4 FILLER_72_919 ();
 fill_1 FILLER_72_923 ();
 fill_2 FILLER_72_925 ();
 fill_4 FILLER_72_936 ();
 fill_2 FILLER_72_940 ();
 fill_1 FILLER_72_942 ();
 fill_2 FILLER_72_949 ();
 fill_1 FILLER_72_951 ();
 fill_2 FILLER_72_956 ();
 fill_1 FILLER_72_979 ();
 fill_8 FILLER_72_996 ();
 fill_2 FILLER_72_1004 ();
 fill_1 FILLER_72_1006 ();
 fill_8 FILLER_72_1025 ();
 fill_1 FILLER_72_1037 ();
 fill_2 FILLER_73_87 ();
 fill_1 FILLER_73_89 ();
 fill_4 FILLER_73_105 ();
 fill_2 FILLER_73_134 ();
 fill_2 FILLER_73_161 ();
 fill_1 FILLER_73_169 ();
 fill_1 FILLER_73_177 ();
 fill_2 FILLER_73_222 ();
 fill_4 FILLER_73_225 ();
 fill_2 FILLER_73_234 ();
 fill_8 FILLER_73_270 ();
 fill_2 FILLER_73_278 ();
 fill_2 FILLER_73_281 ();
 fill_1 FILLER_73_283 ();
 fill_4 FILLER_73_307 ();
 fill_2 FILLER_73_334 ();
 fill_2 FILLER_73_350 ();
 fill_1 FILLER_73_352 ();
 fill_8 FILLER_73_360 ();
 fill_4 FILLER_73_376 ();
 fill_2 FILLER_73_380 ();
 fill_2 FILLER_73_389 ();
 fill_1 FILLER_73_391 ();
 fill_4 FILLER_73_400 ();
 fill_1 FILLER_73_407 ();
 fill_1 FILLER_73_447 ();
 fill_1 FILLER_73_505 ();
 fill_2 FILLER_73_539 ();
 fill_1 FILLER_73_541 ();
 fill_4 FILLER_73_561 ();
 fill_2 FILLER_73_575 ();
 fill_2 FILLER_73_601 ();
 fill_2 FILLER_73_606 ();
 fill_1 FILLER_73_608 ();
 fill_1 FILLER_73_634 ();
 decap_12 FILLER_73_642 ();
 decap_12 FILLER_73_654 ();
 fill_4 FILLER_73_666 ();
 fill_2 FILLER_73_670 ();
 fill_4 FILLER_73_673 ();
 fill_2 FILLER_73_677 ();
 fill_1 FILLER_73_679 ();
 fill_1 FILLER_73_687 ();
 fill_2 FILLER_73_735 ();
 fill_1 FILLER_73_744 ();
 fill_1 FILLER_73_762 ();
 fill_4 FILLER_73_779 ();
 fill_1 FILLER_73_783 ();
 fill_4 FILLER_73_844 ();
 fill_1 FILLER_73_863 ();
 fill_2 FILLER_73_894 ();
 fill_8 FILLER_73_944 ();
 fill_1 FILLER_73_973 ();
 decap_12 FILLER_73_980 ();
 fill_8 FILLER_73_992 ();
 fill_2 FILLER_73_1000 ();
 fill_8 FILLER_73_1029 ();
 fill_1 FILLER_73_1037 ();
 fill_2 FILLER_74_3 ();
 fill_2 FILLER_74_36 ();
 fill_2 FILLER_74_63 ();
 fill_1 FILLER_74_73 ();
 fill_1 FILLER_74_83 ();
 fill_2 FILLER_74_93 ();
 decap_12 FILLER_74_103 ();
 fill_2 FILLER_74_115 ();
 fill_1 FILLER_74_145 ();
 fill_2 FILLER_74_182 ();
 fill_1 FILLER_74_191 ();
 fill_2 FILLER_74_197 ();
 fill_2 FILLER_74_206 ();
 fill_1 FILLER_74_208 ();
 fill_2 FILLER_74_216 ();
 fill_1 FILLER_74_239 ();
 fill_2 FILLER_74_249 ();
 fill_1 FILLER_74_251 ();
 fill_4 FILLER_74_253 ();
 fill_1 FILLER_74_275 ();
 fill_1 FILLER_74_288 ();
 fill_1 FILLER_74_294 ();
 fill_2 FILLER_74_344 ();
 fill_1 FILLER_74_346 ();
 fill_1 FILLER_74_365 ();
 fill_1 FILLER_74_373 ();
 fill_2 FILLER_74_404 ();
 fill_1 FILLER_74_406 ();
 fill_2 FILLER_74_418 ();
 fill_4 FILLER_74_437 ();
 fill_2 FILLER_74_449 ();
 fill_1 FILLER_74_461 ();
 fill_1 FILLER_74_475 ();
 decap_12 FILLER_74_497 ();
 fill_8 FILLER_74_522 ();
 fill_2 FILLER_74_530 ();
 fill_2 FILLER_74_539 ();
 fill_1 FILLER_74_541 ();
 fill_4 FILLER_74_554 ();
 fill_1 FILLER_74_558 ();
 decap_12 FILLER_74_573 ();
 fill_2 FILLER_74_585 ();
 fill_1 FILLER_74_587 ();
 fill_8 FILLER_74_589 ();
 fill_1 FILLER_74_597 ();
 decap_12 FILLER_74_605 ();
 fill_4 FILLER_74_617 ();
 fill_2 FILLER_74_621 ();
 fill_1 FILLER_74_623 ();
 fill_2 FILLER_74_631 ();
 fill_1 FILLER_74_633 ();
 fill_2 FILLER_74_661 ();
 fill_4 FILLER_74_693 ();
 fill_1 FILLER_74_724 ();
 decap_12 FILLER_74_771 ();
 fill_4 FILLER_74_783 ();
 decap_12 FILLER_74_791 ();
 fill_8 FILLER_74_803 ();
 fill_1 FILLER_74_811 ();
 decap_12 FILLER_74_828 ();
 fill_4 FILLER_74_840 ();
 fill_2 FILLER_74_844 ();
 fill_2 FILLER_74_866 ();
 fill_4 FILLER_74_889 ();
 fill_2 FILLER_74_893 ();
 fill_1 FILLER_74_895 ();
 fill_8 FILLER_74_902 ();
 fill_1 FILLER_74_910 ();
 fill_8 FILLER_74_914 ();
 fill_2 FILLER_74_922 ();
 decap_12 FILLER_74_945 ();
 fill_2 FILLER_74_957 ();
 fill_2 FILLER_74_965 ();
 fill_1 FILLER_74_967 ();
 fill_8 FILLER_74_971 ();
 fill_1 FILLER_74_979 ();
 decap_12 FILLER_74_981 ();
 decap_12 FILLER_74_993 ();
 decap_12 FILLER_74_1005 ();
 decap_12 FILLER_74_1017 ();
 fill_4 FILLER_74_1029 ();
 fill_2 FILLER_74_1033 ();
 fill_1 FILLER_74_1035 ();
 fill_1 FILLER_74_1037 ();
 fill_2 FILLER_75_57 ();
 fill_2 FILLER_75_78 ();
 fill_8 FILLER_75_102 ();
 fill_2 FILLER_75_110 ();
 fill_4 FILLER_75_120 ();
 fill_2 FILLER_75_124 ();
 fill_4 FILLER_75_130 ();
 fill_2 FILLER_75_134 ();
 fill_4 FILLER_75_144 ();
 fill_1 FILLER_75_159 ();
 fill_1 FILLER_75_181 ();
 fill_1 FILLER_75_199 ();
 fill_2 FILLER_75_207 ();
 fill_2 FILLER_75_222 ();
 fill_2 FILLER_75_231 ();
 fill_2 FILLER_75_239 ();
 fill_1 FILLER_75_241 ();
 fill_2 FILLER_75_253 ();
 fill_1 FILLER_75_255 ();
 fill_2 FILLER_75_261 ();
 fill_2 FILLER_75_277 ();
 fill_1 FILLER_75_279 ();
 fill_1 FILLER_75_306 ();
 fill_2 FILLER_75_349 ();
 fill_4 FILLER_75_363 ();
 fill_2 FILLER_75_367 ();
 fill_2 FILLER_75_377 ();
 fill_1 FILLER_75_379 ();
 fill_2 FILLER_75_393 ();
 fill_8 FILLER_75_415 ();
 fill_2 FILLER_75_432 ();
 fill_1 FILLER_75_434 ();
 fill_1 FILLER_75_458 ();
 fill_2 FILLER_75_472 ();
 fill_1 FILLER_75_474 ();
 fill_2 FILLER_75_485 ();
 fill_1 FILLER_75_496 ();
 fill_4 FILLER_75_512 ();
 fill_2 FILLER_75_516 ();
 fill_1 FILLER_75_518 ();
 fill_8 FILLER_75_535 ();
 fill_1 FILLER_75_552 ();
 fill_1 FILLER_75_559 ();
 decap_12 FILLER_75_561 ();
 fill_2 FILLER_75_573 ();
 fill_8 FILLER_75_589 ();
 fill_4 FILLER_75_604 ();
 decap_12 FILLER_75_617 ();
 fill_1 FILLER_75_629 ();
 decap_12 FILLER_75_636 ();
 fill_1 FILLER_75_648 ();
 fill_4 FILLER_75_666 ();
 fill_2 FILLER_75_670 ();
 fill_4 FILLER_75_686 ();
 fill_1 FILLER_75_690 ();
 fill_2 FILLER_75_719 ();
 fill_1 FILLER_75_721 ();
 fill_1 FILLER_75_729 ();
 fill_2 FILLER_75_763 ();
 fill_4 FILLER_75_778 ();
 fill_2 FILLER_75_782 ();
 decap_12 FILLER_75_805 ();
 decap_12 FILLER_75_817 ();
 fill_8 FILLER_75_829 ();
 fill_2 FILLER_75_837 ();
 fill_1 FILLER_75_839 ();
 decap_12 FILLER_75_841 ();
 decap_12 FILLER_75_853 ();
 decap_12 FILLER_75_865 ();
 decap_12 FILLER_75_877 ();
 fill_4 FILLER_75_889 ();
 fill_2 FILLER_75_893 ();
 fill_1 FILLER_75_895 ();
 decap_12 FILLER_75_897 ();
 decap_12 FILLER_75_909 ();
 decap_12 FILLER_75_921 ();
 decap_12 FILLER_75_933 ();
 fill_4 FILLER_75_945 ();
 fill_2 FILLER_75_949 ();
 fill_1 FILLER_75_951 ();
 decap_12 FILLER_75_953 ();
 decap_12 FILLER_75_965 ();
 decap_12 FILLER_75_977 ();
 decap_12 FILLER_75_989 ();
 fill_4 FILLER_75_1001 ();
 fill_2 FILLER_75_1005 ();
 fill_1 FILLER_75_1007 ();
 decap_12 FILLER_75_1009 ();
 decap_12 FILLER_75_1021 ();
 fill_4 FILLER_75_1033 ();
 fill_1 FILLER_75_1037 ();
 fill_2 FILLER_76_3 ();
 fill_1 FILLER_76_5 ();
 fill_1 FILLER_76_13 ();
 fill_1 FILLER_76_27 ();
 decap_12 FILLER_76_29 ();
 fill_1 FILLER_76_52 ();
 fill_4 FILLER_76_61 ();
 fill_4 FILLER_76_73 ();
 fill_2 FILLER_76_81 ();
 fill_1 FILLER_76_83 ();
 fill_4 FILLER_76_106 ();
 fill_2 FILLER_76_110 ();
 fill_2 FILLER_76_119 ();
 fill_1 FILLER_76_121 ();
 fill_2 FILLER_76_130 ();
 fill_2 FILLER_76_145 ();
 fill_1 FILLER_76_147 ();
 fill_1 FILLER_76_189 ();
 fill_2 FILLER_76_204 ();
 fill_1 FILLER_76_206 ();
 fill_2 FILLER_76_213 ();
 fill_1 FILLER_76_215 ();
 fill_2 FILLER_76_231 ();
 fill_8 FILLER_76_275 ();
 fill_2 FILLER_76_283 ();
 fill_1 FILLER_76_296 ();
 fill_2 FILLER_76_306 ();
 fill_4 FILLER_76_358 ();
 fill_2 FILLER_76_362 ();
 fill_4 FILLER_76_372 ();
 fill_4 FILLER_76_380 ();
 fill_1 FILLER_76_384 ();
 fill_8 FILLER_76_395 ();
 fill_2 FILLER_76_403 ();
 fill_1 FILLER_76_405 ();
 fill_2 FILLER_76_425 ();
 fill_1 FILLER_76_427 ();
 fill_4 FILLER_76_485 ();
 fill_1 FILLER_76_489 ();
 fill_2 FILLER_76_504 ();
 fill_1 FILLER_76_525 ();
 fill_4 FILLER_76_533 ();
 fill_4 FILLER_76_550 ();
 fill_2 FILLER_76_554 ();
 fill_1 FILLER_76_556 ();
 decap_12 FILLER_76_574 ();
 fill_2 FILLER_76_586 ();
 fill_1 FILLER_76_589 ();
 decap_12 FILLER_76_597 ();
 fill_4 FILLER_76_609 ();
 fill_2 FILLER_76_613 ();
 fill_2 FILLER_76_642 ();
 fill_2 FILLER_76_656 ();
 fill_1 FILLER_76_668 ();
 fill_1 FILLER_76_757 ();
 fill_4 FILLER_76_807 ();
 fill_1 FILLER_76_811 ();
 decap_12 FILLER_76_813 ();
 decap_12 FILLER_76_825 ();
 decap_12 FILLER_76_837 ();
 decap_12 FILLER_76_849 ();
 fill_4 FILLER_76_861 ();
 fill_2 FILLER_76_865 ();
 fill_1 FILLER_76_867 ();
 decap_12 FILLER_76_869 ();
 decap_12 FILLER_76_881 ();
 decap_12 FILLER_76_893 ();
 decap_12 FILLER_76_905 ();
 fill_4 FILLER_76_917 ();
 fill_2 FILLER_76_921 ();
 fill_1 FILLER_76_923 ();
 decap_12 FILLER_76_925 ();
 decap_12 FILLER_76_937 ();
 decap_12 FILLER_76_949 ();
 decap_12 FILLER_76_961 ();
 fill_4 FILLER_76_973 ();
 fill_2 FILLER_76_977 ();
 fill_1 FILLER_76_979 ();
 decap_12 FILLER_76_981 ();
 decap_12 FILLER_76_993 ();
 decap_12 FILLER_76_1005 ();
 decap_12 FILLER_76_1017 ();
 fill_4 FILLER_76_1029 ();
 fill_2 FILLER_76_1033 ();
 fill_1 FILLER_76_1035 ();
 fill_1 FILLER_76_1037 ();
 fill_2 FILLER_77_20 ();
 fill_1 FILLER_77_22 ();
 fill_2 FILLER_77_39 ();
 fill_2 FILLER_77_57 ();
 fill_2 FILLER_77_85 ();
 fill_1 FILLER_77_87 ();
 decap_12 FILLER_77_96 ();
 fill_4 FILLER_77_108 ();
 fill_8 FILLER_77_121 ();
 fill_1 FILLER_77_129 ();
 fill_4 FILLER_77_138 ();
 fill_2 FILLER_77_142 ();
 fill_1 FILLER_77_164 ();
 fill_1 FILLER_77_179 ();
 fill_2 FILLER_77_198 ();
 fill_4 FILLER_77_220 ();
 fill_1 FILLER_77_237 ();
 fill_1 FILLER_77_279 ();
 fill_4 FILLER_77_296 ();
 fill_1 FILLER_77_300 ();
 fill_1 FILLER_77_311 ();
 fill_1 FILLER_77_323 ();
 fill_2 FILLER_77_334 ();
 fill_1 FILLER_77_345 ();
 fill_2 FILLER_77_409 ();
 fill_2 FILLER_77_414 ();
 fill_1 FILLER_77_416 ();
 fill_1 FILLER_77_433 ();
 fill_1 FILLER_77_447 ();
 fill_1 FILLER_77_496 ();
 fill_2 FILLER_77_501 ();
 fill_1 FILLER_77_503 ();
 fill_2 FILLER_77_508 ();
 fill_1 FILLER_77_510 ();
 fill_2 FILLER_77_521 ();
 fill_1 FILLER_77_523 ();
 fill_1 FILLER_77_541 ();
 fill_4 FILLER_77_555 ();
 fill_1 FILLER_77_559 ();
 fill_2 FILLER_77_582 ();
 fill_1 FILLER_77_584 ();
 fill_2 FILLER_77_599 ();
 fill_1 FILLER_77_601 ();
 fill_1 FILLER_77_605 ();
 fill_4 FILLER_77_610 ();
 fill_2 FILLER_77_614 ();
 fill_8 FILLER_77_634 ();
 fill_1 FILLER_77_642 ();
 fill_8 FILLER_77_673 ();
 fill_2 FILLER_77_681 ();
 fill_1 FILLER_77_683 ();
 fill_1 FILLER_77_732 ();
 fill_1 FILLER_77_744 ();
 fill_2 FILLER_77_771 ();
 fill_2 FILLER_77_782 ();
 decap_12 FILLER_77_823 ();
 fill_4 FILLER_77_835 ();
 fill_1 FILLER_77_839 ();
 decap_12 FILLER_77_841 ();
 decap_12 FILLER_77_853 ();
 decap_12 FILLER_77_865 ();
 decap_12 FILLER_77_877 ();
 fill_4 FILLER_77_889 ();
 fill_2 FILLER_77_893 ();
 fill_1 FILLER_77_895 ();
 decap_12 FILLER_77_897 ();
 decap_12 FILLER_77_909 ();
 decap_12 FILLER_77_921 ();
 decap_12 FILLER_77_933 ();
 fill_4 FILLER_77_945 ();
 fill_2 FILLER_77_949 ();
 fill_1 FILLER_77_951 ();
 decap_12 FILLER_77_953 ();
 decap_12 FILLER_77_965 ();
 decap_12 FILLER_77_977 ();
 decap_12 FILLER_77_989 ();
 fill_4 FILLER_77_1001 ();
 fill_2 FILLER_77_1005 ();
 fill_1 FILLER_77_1007 ();
 decap_12 FILLER_77_1009 ();
 decap_12 FILLER_77_1021 ();
 fill_4 FILLER_77_1033 ();
 fill_1 FILLER_77_1037 ();
 fill_2 FILLER_78_3 ();
 fill_2 FILLER_78_16 ();
 fill_4 FILLER_78_62 ();
 fill_2 FILLER_78_66 ();
 fill_4 FILLER_78_79 ();
 fill_1 FILLER_78_83 ();
 fill_4 FILLER_78_85 ();
 fill_2 FILLER_78_89 ();
 fill_1 FILLER_78_104 ();
 fill_4 FILLER_78_122 ();
 fill_1 FILLER_78_126 ();
 fill_4 FILLER_78_135 ();
 fill_1 FILLER_78_139 ();
 fill_8 FILLER_78_141 ();
 fill_2 FILLER_78_149 ();
 fill_1 FILLER_78_151 ();
 fill_4 FILLER_78_160 ();
 fill_2 FILLER_78_188 ();
 fill_2 FILLER_78_214 ();
 fill_8 FILLER_78_225 ();
 fill_1 FILLER_78_233 ();
 fill_2 FILLER_78_250 ();
 fill_1 FILLER_78_257 ();
 fill_1 FILLER_78_275 ();
 fill_4 FILLER_78_312 ();
 fill_2 FILLER_78_316 ();
 fill_2 FILLER_78_335 ();
 fill_4 FILLER_78_342 ();
 fill_2 FILLER_78_346 ();
 fill_1 FILLER_78_348 ();
 fill_8 FILLER_78_354 ();
 fill_2 FILLER_78_362 ();
 fill_4 FILLER_78_369 ();
 fill_2 FILLER_78_373 ();
 fill_1 FILLER_78_375 ();
 fill_8 FILLER_78_389 ();
 fill_1 FILLER_78_397 ();
 fill_8 FILLER_78_412 ();
 fill_2 FILLER_78_421 ();
 fill_1 FILLER_78_439 ();
 fill_2 FILLER_78_533 ();
 fill_8 FILLER_78_561 ();
 fill_4 FILLER_78_582 ();
 fill_2 FILLER_78_586 ();
 fill_2 FILLER_78_589 ();
 fill_1 FILLER_78_591 ();
 fill_2 FILLER_78_599 ();
 fill_2 FILLER_78_613 ();
 fill_1 FILLER_78_615 ();
 fill_2 FILLER_78_629 ();
 fill_1 FILLER_78_631 ();
 fill_2 FILLER_78_642 ();
 fill_4 FILLER_78_652 ();
 fill_1 FILLER_78_707 ();
 fill_4 FILLER_78_724 ();
 fill_1 FILLER_78_728 ();
 fill_2 FILLER_78_740 ();
 fill_4 FILLER_78_806 ();
 fill_2 FILLER_78_810 ();
 fill_2 FILLER_78_813 ();
 fill_1 FILLER_78_815 ();
 decap_12 FILLER_78_825 ();
 decap_12 FILLER_78_837 ();
 decap_12 FILLER_78_849 ();
 fill_4 FILLER_78_861 ();
 fill_2 FILLER_78_865 ();
 fill_1 FILLER_78_867 ();
 decap_12 FILLER_78_869 ();
 decap_12 FILLER_78_881 ();
 decap_12 FILLER_78_893 ();
 decap_12 FILLER_78_905 ();
 fill_4 FILLER_78_917 ();
 fill_2 FILLER_78_921 ();
 fill_1 FILLER_78_923 ();
 decap_12 FILLER_78_925 ();
 decap_12 FILLER_78_937 ();
 decap_12 FILLER_78_949 ();
 decap_12 FILLER_78_961 ();
 fill_4 FILLER_78_973 ();
 fill_2 FILLER_78_977 ();
 fill_1 FILLER_78_979 ();
 decap_12 FILLER_78_981 ();
 decap_12 FILLER_78_993 ();
 decap_12 FILLER_78_1005 ();
 decap_12 FILLER_78_1017 ();
 fill_4 FILLER_78_1029 ();
 fill_2 FILLER_78_1033 ();
 fill_1 FILLER_78_1035 ();
 fill_1 FILLER_78_1037 ();
 fill_4 FILLER_79_3 ();
 fill_2 FILLER_79_7 ();
 fill_1 FILLER_79_26 ();
 fill_2 FILLER_79_54 ();
 fill_2 FILLER_79_57 ();
 fill_2 FILLER_79_67 ();
 fill_4 FILLER_79_105 ();
 fill_2 FILLER_79_109 ();
 fill_1 FILLER_79_111 ();
 fill_8 FILLER_79_113 ();
 fill_2 FILLER_79_121 ();
 fill_1 FILLER_79_123 ();
 fill_2 FILLER_79_141 ();
 fill_8 FILLER_79_157 ();
 fill_2 FILLER_79_165 ();
 fill_1 FILLER_79_167 ();
 fill_2 FILLER_79_172 ();
 fill_1 FILLER_79_174 ();
 fill_2 FILLER_79_181 ();
 fill_1 FILLER_79_202 ();
 fill_4 FILLER_79_211 ();
 fill_1 FILLER_79_215 ();
 fill_1 FILLER_79_225 ();
 fill_4 FILLER_79_234 ();
 fill_1 FILLER_79_238 ();
 fill_1 FILLER_79_253 ();
 fill_1 FILLER_79_259 ();
 fill_2 FILLER_79_265 ();
 fill_4 FILLER_79_273 ();
 fill_2 FILLER_79_277 ();
 fill_1 FILLER_79_279 ();
 decap_12 FILLER_79_281 ();
 fill_4 FILLER_79_293 ();
 fill_1 FILLER_79_313 ();
 fill_4 FILLER_79_319 ();
 fill_2 FILLER_79_323 ();
 fill_1 FILLER_79_325 ();
 fill_4 FILLER_79_331 ();
 fill_1 FILLER_79_335 ();
 fill_4 FILLER_79_337 ();
 fill_4 FILLER_79_357 ();
 fill_1 FILLER_79_361 ();
 fill_4 FILLER_79_370 ();
 fill_2 FILLER_79_374 ();
 fill_2 FILLER_79_400 ();
 fill_1 FILLER_79_402 ();
 fill_8 FILLER_79_417 ();
 fill_1 FILLER_79_425 ();
 fill_2 FILLER_79_438 ();
 fill_2 FILLER_79_446 ();
 fill_1 FILLER_79_453 ();
 fill_1 FILLER_79_463 ();
 fill_4 FILLER_79_475 ();
 fill_2 FILLER_79_495 ();
 fill_1 FILLER_79_503 ();
 fill_2 FILLER_79_505 ();
 fill_2 FILLER_79_532 ();
 fill_4 FILLER_79_537 ();
 fill_2 FILLER_79_561 ();
 fill_4 FILLER_79_592 ();
 decap_12 FILLER_79_603 ();
 fill_1 FILLER_79_615 ();
 fill_2 FILLER_79_624 ();
 fill_4 FILLER_79_639 ();
 fill_1 FILLER_79_643 ();
 fill_2 FILLER_79_660 ();
 fill_1 FILLER_79_673 ();
 fill_1 FILLER_79_735 ();
 fill_1 FILLER_79_776 ();
 fill_1 FILLER_79_785 ();
 fill_4 FILLER_79_833 ();
 fill_2 FILLER_79_837 ();
 fill_1 FILLER_79_839 ();
 decap_12 FILLER_79_841 ();
 decap_12 FILLER_79_853 ();
 decap_12 FILLER_79_865 ();
 decap_12 FILLER_79_877 ();
 fill_4 FILLER_79_889 ();
 fill_2 FILLER_79_893 ();
 fill_1 FILLER_79_895 ();
 decap_12 FILLER_79_897 ();
 decap_12 FILLER_79_909 ();
 decap_12 FILLER_79_921 ();
 decap_12 FILLER_79_933 ();
 fill_4 FILLER_79_945 ();
 fill_2 FILLER_79_949 ();
 fill_1 FILLER_79_951 ();
 decap_12 FILLER_79_953 ();
 decap_12 FILLER_79_965 ();
 decap_12 FILLER_79_977 ();
 decap_12 FILLER_79_989 ();
 fill_4 FILLER_79_1001 ();
 fill_2 FILLER_79_1005 ();
 fill_1 FILLER_79_1007 ();
 decap_12 FILLER_79_1009 ();
 decap_12 FILLER_79_1021 ();
 fill_4 FILLER_79_1033 ();
 fill_1 FILLER_79_1037 ();
 fill_2 FILLER_80_19 ();
 fill_1 FILLER_80_79 ();
 fill_1 FILLER_80_83 ();
 decap_12 FILLER_80_93 ();
 decap_12 FILLER_80_105 ();
 fill_4 FILLER_80_117 ();
 fill_1 FILLER_80_121 ();
 fill_4 FILLER_80_130 ();
 fill_2 FILLER_80_134 ();
 fill_4 FILLER_80_168 ();
 fill_2 FILLER_80_172 ();
 fill_8 FILLER_80_186 ();
 fill_2 FILLER_80_194 ();
 fill_4 FILLER_80_212 ();
 fill_2 FILLER_80_216 ();
 decap_12 FILLER_80_225 ();
 fill_2 FILLER_80_237 ();
 fill_1 FILLER_80_239 ();
 fill_4 FILLER_80_248 ();
 fill_4 FILLER_80_253 ();
 fill_8 FILLER_80_265 ();
 fill_2 FILLER_80_278 ();
 decap_12 FILLER_80_288 ();
 fill_8 FILLER_80_300 ();
 decap_12 FILLER_80_309 ();
 fill_8 FILLER_80_328 ();
 decap_12 FILLER_80_343 ();
 fill_2 FILLER_80_355 ();
 fill_2 FILLER_80_365 ();
 fill_4 FILLER_80_381 ();
 fill_1 FILLER_80_385 ();
 decap_12 FILLER_80_394 ();
 fill_8 FILLER_80_406 ();
 fill_2 FILLER_80_414 ();
 fill_1 FILLER_80_416 ();
 fill_1 FILLER_80_449 ();
 fill_4 FILLER_80_489 ();
 fill_1 FILLER_80_493 ();
 fill_1 FILLER_80_531 ();
 fill_2 FILLER_80_533 ();
 fill_1 FILLER_80_543 ();
 fill_2 FILLER_80_558 ();
 fill_1 FILLER_80_569 ();
 fill_8 FILLER_80_579 ();
 fill_1 FILLER_80_587 ();
 fill_1 FILLER_80_606 ();
 fill_4 FILLER_80_621 ();
 decap_12 FILLER_80_629 ();
 fill_2 FILLER_80_641 ();
 fill_1 FILLER_80_643 ();
 fill_4 FILLER_80_645 ();
 fill_2 FILLER_80_793 ();
 fill_2 FILLER_80_813 ();
 fill_1 FILLER_80_815 ();
 decap_12 FILLER_80_837 ();
 decap_12 FILLER_80_849 ();
 fill_4 FILLER_80_861 ();
 fill_2 FILLER_80_865 ();
 fill_1 FILLER_80_867 ();
 decap_12 FILLER_80_869 ();
 decap_12 FILLER_80_881 ();
 decap_12 FILLER_80_893 ();
 decap_12 FILLER_80_905 ();
 fill_4 FILLER_80_917 ();
 fill_2 FILLER_80_921 ();
 fill_1 FILLER_80_923 ();
 decap_12 FILLER_80_925 ();
 decap_12 FILLER_80_937 ();
 decap_12 FILLER_80_949 ();
 decap_12 FILLER_80_961 ();
 fill_4 FILLER_80_973 ();
 fill_2 FILLER_80_977 ();
 fill_1 FILLER_80_979 ();
 decap_12 FILLER_80_981 ();
 decap_12 FILLER_80_993 ();
 decap_12 FILLER_80_1005 ();
 decap_12 FILLER_80_1017 ();
 fill_4 FILLER_80_1029 ();
 fill_2 FILLER_80_1033 ();
 fill_1 FILLER_80_1035 ();
 fill_1 FILLER_80_1037 ();
 fill_8 FILLER_81_3 ();
 fill_2 FILLER_81_22 ();
 fill_8 FILLER_81_31 ();
 fill_1 FILLER_81_55 ();
 fill_4 FILLER_81_100 ();
 fill_1 FILLER_81_104 ();
 fill_1 FILLER_81_128 ();
 fill_1 FILLER_81_137 ();
 fill_4 FILLER_81_169 ();
 fill_1 FILLER_81_173 ();
 fill_4 FILLER_81_182 ();
 fill_1 FILLER_81_186 ();
 fill_1 FILLER_81_208 ();
 fill_4 FILLER_81_217 ();
 fill_2 FILLER_81_221 ();
 fill_1 FILLER_81_223 ();
 decap_12 FILLER_81_233 ();
 fill_8 FILLER_81_245 ();
 fill_2 FILLER_81_253 ();
 decap_12 FILLER_81_263 ();
 fill_4 FILLER_81_275 ();
 fill_1 FILLER_81_279 ();
 fill_8 FILLER_81_281 ();
 fill_2 FILLER_81_289 ();
 fill_4 FILLER_81_299 ();
 fill_2 FILLER_81_303 ();
 fill_1 FILLER_81_305 ();
 fill_4 FILLER_81_322 ();
 fill_2 FILLER_81_326 ();
 fill_1 FILLER_81_337 ();
 fill_4 FILLER_81_345 ();
 fill_1 FILLER_81_349 ();
 fill_1 FILLER_81_364 ();
 fill_2 FILLER_81_369 ();
 fill_1 FILLER_81_371 ();
 fill_4 FILLER_81_386 ();
 fill_2 FILLER_81_390 ();
 fill_2 FILLER_81_393 ();
 fill_1 FILLER_81_395 ();
 fill_2 FILLER_81_403 ();
 fill_1 FILLER_81_405 ();
 decap_12 FILLER_81_413 ();
 fill_2 FILLER_81_425 ();
 fill_1 FILLER_81_427 ();
 fill_1 FILLER_81_464 ();
 fill_4 FILLER_81_499 ();
 fill_1 FILLER_81_503 ();
 fill_1 FILLER_81_517 ();
 fill_4 FILLER_81_534 ();
 fill_1 FILLER_81_538 ();
 fill_1 FILLER_81_542 ();
 fill_2 FILLER_81_558 ();
 fill_2 FILLER_81_585 ();
 fill_4 FILLER_81_650 ();
 fill_1 FILLER_81_654 ();
 fill_1 FILLER_81_680 ();
 fill_1 FILLER_81_755 ();
 fill_2 FILLER_81_777 ();
 fill_1 FILLER_81_779 ();
 fill_4 FILLER_81_835 ();
 fill_1 FILLER_81_839 ();
 decap_12 FILLER_81_841 ();
 decap_12 FILLER_81_853 ();
 decap_12 FILLER_81_865 ();
 decap_12 FILLER_81_877 ();
 fill_4 FILLER_81_889 ();
 fill_2 FILLER_81_893 ();
 fill_1 FILLER_81_895 ();
 decap_12 FILLER_81_897 ();
 decap_12 FILLER_81_909 ();
 decap_12 FILLER_81_921 ();
 decap_12 FILLER_81_933 ();
 fill_4 FILLER_81_945 ();
 fill_2 FILLER_81_949 ();
 fill_1 FILLER_81_951 ();
 decap_12 FILLER_81_953 ();
 decap_12 FILLER_81_965 ();
 decap_12 FILLER_81_977 ();
 decap_12 FILLER_81_989 ();
 fill_4 FILLER_81_1001 ();
 fill_2 FILLER_81_1005 ();
 fill_1 FILLER_81_1007 ();
 decap_12 FILLER_81_1009 ();
 decap_12 FILLER_81_1021 ();
 fill_1 FILLER_81_1033 ();
 fill_2 FILLER_82_3 ();
 fill_1 FILLER_82_5 ();
 fill_4 FILLER_82_24 ();
 fill_2 FILLER_82_54 ();
 fill_1 FILLER_82_56 ();
 fill_2 FILLER_82_82 ();
 fill_4 FILLER_82_85 ();
 fill_4 FILLER_82_166 ();
 fill_2 FILLER_82_170 ();
 fill_8 FILLER_82_176 ();
 fill_1 FILLER_82_184 ();
 fill_4 FILLER_82_192 ();
 fill_4 FILLER_82_211 ();
 fill_2 FILLER_82_215 ();
 fill_8 FILLER_82_242 ();
 fill_2 FILLER_82_250 ();
 fill_2 FILLER_82_253 ();
 fill_1 FILLER_82_255 ();
 fill_8 FILLER_82_263 ();
 decap_12 FILLER_82_293 ();
 fill_2 FILLER_82_305 ();
 fill_1 FILLER_82_307 ();
 decap_12 FILLER_82_309 ();
 fill_8 FILLER_82_321 ();
 fill_1 FILLER_82_352 ();
 fill_2 FILLER_82_361 ();
 fill_1 FILLER_82_363 ();
 fill_2 FILLER_82_365 ();
 fill_1 FILLER_82_367 ();
 fill_2 FILLER_82_373 ();
 fill_1 FILLER_82_375 ();
 fill_2 FILLER_82_424 ();
 fill_1 FILLER_82_426 ();
 fill_1 FILLER_82_475 ();
 fill_2 FILLER_82_477 ();
 fill_1 FILLER_82_523 ();
 fill_4 FILLER_82_527 ();
 fill_1 FILLER_82_531 ();
 fill_2 FILLER_82_533 ();
 fill_2 FILLER_82_538 ();
 fill_1 FILLER_82_540 ();
 fill_1 FILLER_82_587 ();
 decap_12 FILLER_82_604 ();
 decap_12 FILLER_82_616 ();
 decap_12 FILLER_82_628 ();
 fill_4 FILLER_82_640 ();
 fill_1 FILLER_82_645 ();
 fill_8 FILLER_82_649 ();
 fill_2 FILLER_82_657 ();
 fill_1 FILLER_82_659 ();
 fill_2 FILLER_82_706 ();
 fill_2 FILLER_82_715 ();
 fill_2 FILLER_82_725 ();
 fill_4 FILLER_82_750 ();
 fill_2 FILLER_82_754 ();
 fill_2 FILLER_82_799 ();
 fill_1 FILLER_82_801 ();
 fill_1 FILLER_82_811 ();
 decap_12 FILLER_82_840 ();
 decap_12 FILLER_82_852 ();
 fill_4 FILLER_82_864 ();
 decap_12 FILLER_82_869 ();
 decap_12 FILLER_82_881 ();
 decap_12 FILLER_82_893 ();
 decap_12 FILLER_82_905 ();
 fill_4 FILLER_82_917 ();
 fill_2 FILLER_82_921 ();
 fill_1 FILLER_82_923 ();
 decap_12 FILLER_82_925 ();
 decap_12 FILLER_82_937 ();
 decap_12 FILLER_82_949 ();
 decap_12 FILLER_82_961 ();
 fill_4 FILLER_82_973 ();
 fill_2 FILLER_82_977 ();
 fill_1 FILLER_82_979 ();
 decap_12 FILLER_82_981 ();
 decap_12 FILLER_82_993 ();
 decap_12 FILLER_82_1005 ();
 decap_12 FILLER_82_1017 ();
 fill_4 FILLER_82_1029 ();
 fill_2 FILLER_82_1033 ();
 fill_1 FILLER_82_1035 ();
 fill_1 FILLER_82_1037 ();
 fill_4 FILLER_83_41 ();
 fill_1 FILLER_83_45 ();
 fill_2 FILLER_83_54 ();
 fill_4 FILLER_83_57 ();
 fill_4 FILLER_83_78 ();
 fill_4 FILLER_83_99 ();
 fill_2 FILLER_83_103 ();
 fill_2 FILLER_83_146 ();
 fill_1 FILLER_83_169 ();
 fill_8 FILLER_83_186 ();
 fill_4 FILLER_83_213 ();
 fill_2 FILLER_83_233 ();
 fill_4 FILLER_83_250 ();
 fill_2 FILLER_83_254 ();
 fill_4 FILLER_83_263 ();
 fill_2 FILLER_83_291 ();
 fill_1 FILLER_83_293 ();
 fill_4 FILLER_83_302 ();
 fill_2 FILLER_83_315 ();
 fill_1 FILLER_83_325 ();
 fill_2 FILLER_83_334 ();
 fill_8 FILLER_83_344 ();
 fill_4 FILLER_83_359 ();
 fill_2 FILLER_83_363 ();
 fill_2 FILLER_83_379 ();
 fill_1 FILLER_83_381 ();
 fill_4 FILLER_83_406 ();
 fill_2 FILLER_83_413 ();
 fill_2 FILLER_83_441 ();
 fill_1 FILLER_83_443 ();
 fill_1 FILLER_83_447 ();
 fill_4 FILLER_83_459 ();
 fill_2 FILLER_83_463 ();
 fill_8 FILLER_83_477 ();
 fill_1 FILLER_83_485 ();
 fill_2 FILLER_83_505 ();
 fill_1 FILLER_83_507 ();
 fill_2 FILLER_83_548 ();
 fill_1 FILLER_83_550 ();
 fill_2 FILLER_83_561 ();
 fill_1 FILLER_83_571 ();
 fill_4 FILLER_83_606 ();
 fill_2 FILLER_83_613 ();
 fill_1 FILLER_83_615 ();
 fill_1 FILLER_83_617 ();
 fill_8 FILLER_83_625 ();
 fill_2 FILLER_83_656 ();
 fill_8 FILLER_83_737 ();
 fill_2 FILLER_83_745 ();
 fill_1 FILLER_83_747 ();
 fill_4 FILLER_83_774 ();
 fill_1 FILLER_83_839 ();
 decap_12 FILLER_83_841 ();
 decap_12 FILLER_83_853 ();
 decap_12 FILLER_83_865 ();
 decap_12 FILLER_83_877 ();
 fill_4 FILLER_83_889 ();
 fill_2 FILLER_83_893 ();
 fill_1 FILLER_83_895 ();
 decap_12 FILLER_83_897 ();
 decap_12 FILLER_83_909 ();
 decap_12 FILLER_83_921 ();
 decap_12 FILLER_83_933 ();
 fill_4 FILLER_83_945 ();
 fill_2 FILLER_83_949 ();
 fill_1 FILLER_83_951 ();
 decap_12 FILLER_83_953 ();
 decap_12 FILLER_83_965 ();
 decap_12 FILLER_83_977 ();
 decap_12 FILLER_83_989 ();
 fill_4 FILLER_83_1001 ();
 fill_2 FILLER_83_1005 ();
 fill_1 FILLER_83_1007 ();
 decap_12 FILLER_83_1009 ();
 decap_12 FILLER_83_1021 ();
 fill_4 FILLER_83_1033 ();
 fill_1 FILLER_83_1037 ();
 fill_2 FILLER_84_3 ();
 fill_1 FILLER_84_5 ();
 fill_2 FILLER_84_26 ();
 fill_1 FILLER_84_46 ();
 fill_2 FILLER_84_63 ();
 fill_2 FILLER_84_81 ();
 fill_1 FILLER_84_83 ();
 fill_4 FILLER_84_93 ();
 fill_8 FILLER_84_175 ();
 fill_2 FILLER_84_183 ();
 fill_1 FILLER_84_185 ();
 fill_2 FILLER_84_194 ();
 fill_2 FILLER_84_197 ();
 fill_1 FILLER_84_199 ();
 fill_2 FILLER_84_215 ();
 decap_12 FILLER_84_224 ();
 fill_4 FILLER_84_236 ();
 fill_8 FILLER_84_244 ();
 decap_12 FILLER_84_253 ();
 fill_8 FILLER_84_265 ();
 fill_2 FILLER_84_273 ();
 fill_1 FILLER_84_275 ();
 fill_2 FILLER_84_281 ();
 fill_2 FILLER_84_298 ();
 fill_1 FILLER_84_315 ();
 fill_1 FILLER_84_355 ();
 fill_2 FILLER_84_362 ();
 fill_1 FILLER_84_365 ();
 fill_1 FILLER_84_375 ();
 fill_2 FILLER_84_392 ();
 fill_4 FILLER_84_421 ();
 fill_2 FILLER_84_425 ();
 fill_1 FILLER_84_427 ();
 fill_2 FILLER_84_510 ();
 fill_1 FILLER_84_519 ();
 fill_4 FILLER_84_523 ();
 fill_2 FILLER_84_527 ();
 fill_1 FILLER_84_548 ();
 fill_2 FILLER_84_569 ();
 fill_1 FILLER_84_587 ();
 fill_1 FILLER_84_601 ();
 fill_1 FILLER_84_610 ();
 fill_1 FILLER_84_616 ();
 fill_2 FILLER_84_648 ();
 fill_1 FILLER_84_650 ();
 fill_1 FILLER_84_696 ();
 fill_1 FILLER_84_701 ();
 fill_1 FILLER_84_728 ();
 fill_2 FILLER_84_747 ();
 fill_2 FILLER_84_764 ();
 fill_1 FILLER_84_766 ();
 fill_2 FILLER_84_784 ();
 fill_1 FILLER_84_786 ();
 fill_2 FILLER_84_809 ();
 fill_1 FILLER_84_811 ();
 fill_4 FILLER_84_813 ();
 decap_12 FILLER_84_833 ();
 decap_12 FILLER_84_845 ();
 fill_8 FILLER_84_857 ();
 fill_2 FILLER_84_865 ();
 fill_1 FILLER_84_867 ();
 decap_12 FILLER_84_869 ();
 decap_12 FILLER_84_881 ();
 decap_12 FILLER_84_893 ();
 decap_12 FILLER_84_905 ();
 fill_4 FILLER_84_917 ();
 fill_2 FILLER_84_921 ();
 fill_1 FILLER_84_923 ();
 decap_12 FILLER_84_925 ();
 decap_12 FILLER_84_937 ();
 decap_12 FILLER_84_949 ();
 decap_12 FILLER_84_961 ();
 fill_4 FILLER_84_973 ();
 fill_2 FILLER_84_977 ();
 fill_1 FILLER_84_979 ();
 decap_12 FILLER_84_981 ();
 decap_12 FILLER_84_993 ();
 decap_12 FILLER_84_1005 ();
 decap_12 FILLER_84_1017 ();
 fill_4 FILLER_84_1029 ();
 fill_2 FILLER_84_1033 ();
 fill_1 FILLER_84_1035 ();
 fill_1 FILLER_84_1037 ();
 fill_1 FILLER_85_24 ();
 fill_4 FILLER_85_42 ();
 fill_1 FILLER_85_46 ();
 fill_1 FILLER_85_55 ();
 fill_4 FILLER_85_57 ();
 fill_2 FILLER_85_61 ();
 fill_2 FILLER_85_76 ();
 fill_1 FILLER_85_78 ();
 fill_4 FILLER_85_87 ();
 fill_1 FILLER_85_91 ();
 fill_1 FILLER_85_113 ();
 fill_2 FILLER_85_165 ();
 fill_1 FILLER_85_167 ();
 fill_1 FILLER_85_186 ();
 fill_2 FILLER_85_195 ();
 fill_1 FILLER_85_205 ();
 fill_2 FILLER_85_213 ();
 fill_1 FILLER_85_215 ();
 fill_2 FILLER_85_240 ();
 fill_2 FILLER_85_246 ();
 fill_1 FILLER_85_248 ();
 fill_4 FILLER_85_256 ();
 fill_4 FILLER_85_276 ();
 fill_2 FILLER_85_281 ();
 fill_4 FILLER_85_297 ();
 fill_2 FILLER_85_301 ();
 fill_2 FILLER_85_307 ();
 fill_4 FILLER_85_332 ();
 fill_4 FILLER_85_341 ();
 fill_2 FILLER_85_345 ();
 fill_4 FILLER_85_352 ();
 fill_1 FILLER_85_356 ();
 fill_4 FILLER_85_364 ();
 fill_2 FILLER_85_368 ();
 fill_2 FILLER_85_379 ();
 fill_2 FILLER_85_385 ();
 fill_2 FILLER_85_393 ();
 fill_8 FILLER_85_408 ();
 fill_2 FILLER_85_416 ();
 fill_4 FILLER_85_425 ();
 decap_12 FILLER_85_432 ();
 fill_4 FILLER_85_444 ();
 decap_12 FILLER_85_449 ();
 fill_2 FILLER_85_461 ();
 fill_1 FILLER_85_492 ();
 fill_4 FILLER_85_531 ();
 fill_1 FILLER_85_535 ();
 fill_4 FILLER_85_551 ();
 fill_1 FILLER_85_555 ();
 fill_2 FILLER_85_561 ();
 decap_12 FILLER_85_571 ();
 fill_2 FILLER_85_613 ();
 fill_1 FILLER_85_615 ();
 decap_12 FILLER_85_617 ();
 fill_4 FILLER_85_629 ();
 fill_2 FILLER_85_633 ();
 fill_4 FILLER_85_651 ();
 fill_2 FILLER_85_655 ();
 fill_4 FILLER_85_668 ();
 fill_4 FILLER_85_683 ();
 fill_1 FILLER_85_720 ();
 fill_1 FILLER_85_727 ();
 fill_1 FILLER_85_750 ();
 fill_4 FILLER_85_779 ();
 fill_1 FILLER_85_783 ();
 fill_2 FILLER_85_794 ();
 fill_1 FILLER_85_796 ();
 fill_2 FILLER_85_837 ();
 fill_1 FILLER_85_839 ();
 decap_12 FILLER_85_841 ();
 decap_12 FILLER_85_853 ();
 decap_12 FILLER_85_865 ();
 decap_12 FILLER_85_877 ();
 fill_4 FILLER_85_889 ();
 fill_2 FILLER_85_893 ();
 fill_1 FILLER_85_895 ();
 decap_12 FILLER_85_897 ();
 decap_12 FILLER_85_909 ();
 decap_12 FILLER_85_921 ();
 decap_12 FILLER_85_933 ();
 fill_4 FILLER_85_945 ();
 fill_2 FILLER_85_949 ();
 fill_1 FILLER_85_951 ();
 decap_12 FILLER_85_953 ();
 decap_12 FILLER_85_965 ();
 decap_12 FILLER_85_977 ();
 decap_12 FILLER_85_989 ();
 fill_4 FILLER_85_1001 ();
 fill_2 FILLER_85_1005 ();
 fill_1 FILLER_85_1007 ();
 decap_12 FILLER_85_1009 ();
 decap_12 FILLER_85_1021 ();
 fill_4 FILLER_85_1033 ();
 fill_1 FILLER_85_1037 ();
 fill_4 FILLER_86_3 ();
 fill_2 FILLER_86_7 ();
 fill_1 FILLER_86_16 ();
 fill_4 FILLER_86_22 ();
 fill_2 FILLER_86_26 ();
 fill_2 FILLER_86_51 ();
 fill_1 FILLER_86_53 ();
 fill_2 FILLER_86_81 ();
 fill_1 FILLER_86_83 ();
 fill_4 FILLER_86_104 ();
 fill_2 FILLER_86_108 ();
 fill_1 FILLER_86_110 ();
 decap_12 FILLER_86_128 ();
 fill_4 FILLER_86_148 ();
 fill_1 FILLER_86_152 ();
 fill_2 FILLER_86_193 ();
 fill_1 FILLER_86_195 ();
 fill_2 FILLER_86_197 ();
 fill_1 FILLER_86_199 ();
 fill_4 FILLER_86_210 ();
 fill_2 FILLER_86_299 ();
 fill_4 FILLER_86_309 ();
 fill_1 FILLER_86_313 ();
 fill_4 FILLER_86_353 ();
 fill_1 FILLER_86_385 ();
 fill_1 FILLER_86_391 ();
 fill_2 FILLER_86_395 ();
 fill_1 FILLER_86_401 ();
 fill_2 FILLER_86_417 ();
 fill_1 FILLER_86_419 ();
 fill_1 FILLER_86_432 ();
 fill_2 FILLER_86_452 ();
 fill_1 FILLER_86_465 ();
 fill_8 FILLER_86_536 ();
 fill_2 FILLER_86_549 ();
 fill_1 FILLER_86_551 ();
 fill_1 FILLER_86_561 ();
 fill_1 FILLER_86_587 ();
 fill_4 FILLER_86_589 ();
 fill_1 FILLER_86_593 ();
 decap_12 FILLER_86_597 ();
 fill_8 FILLER_86_614 ();
 fill_2 FILLER_86_622 ();
 fill_1 FILLER_86_624 ();
 fill_4 FILLER_86_631 ();
 fill_1 FILLER_86_635 ();
 fill_1 FILLER_86_658 ();
 fill_2 FILLER_86_668 ();
 fill_1 FILLER_86_670 ();
 fill_2 FILLER_86_680 ();
 fill_1 FILLER_86_682 ();
 fill_4 FILLER_86_695 ();
 fill_1 FILLER_86_699 ();
 fill_4 FILLER_86_701 ();
 fill_1 FILLER_86_734 ();
 fill_8 FILLER_86_794 ();
 fill_1 FILLER_86_811 ();
 fill_1 FILLER_86_819 ();
 decap_12 FILLER_86_847 ();
 fill_8 FILLER_86_859 ();
 fill_1 FILLER_86_867 ();
 decap_12 FILLER_86_869 ();
 decap_12 FILLER_86_881 ();
 decap_12 FILLER_86_893 ();
 decap_12 FILLER_86_905 ();
 fill_4 FILLER_86_917 ();
 fill_2 FILLER_86_921 ();
 fill_1 FILLER_86_923 ();
 decap_12 FILLER_86_925 ();
 decap_12 FILLER_86_937 ();
 decap_12 FILLER_86_949 ();
 decap_12 FILLER_86_961 ();
 fill_4 FILLER_86_973 ();
 fill_2 FILLER_86_977 ();
 fill_1 FILLER_86_979 ();
 decap_12 FILLER_86_981 ();
 decap_12 FILLER_86_993 ();
 decap_12 FILLER_86_1005 ();
 decap_12 FILLER_86_1017 ();
 fill_4 FILLER_86_1029 ();
 fill_2 FILLER_86_1033 ();
 fill_1 FILLER_86_1035 ();
 fill_1 FILLER_86_1037 ();
 fill_4 FILLER_87_32 ();
 fill_2 FILLER_87_36 ();
 fill_4 FILLER_87_50 ();
 fill_2 FILLER_87_54 ();
 fill_2 FILLER_87_84 ();
 fill_1 FILLER_87_92 ();
 fill_4 FILLER_87_100 ();
 fill_2 FILLER_87_104 ();
 fill_1 FILLER_87_106 ();
 fill_1 FILLER_87_113 ();
 fill_2 FILLER_87_166 ();
 decap_12 FILLER_87_178 ();
 fill_4 FILLER_87_205 ();
 fill_2 FILLER_87_222 ();
 fill_4 FILLER_87_225 ();
 fill_2 FILLER_87_245 ();
 fill_2 FILLER_87_253 ();
 fill_1 FILLER_87_255 ();
 fill_2 FILLER_87_277 ();
 fill_1 FILLER_87_279 ();
 fill_1 FILLER_87_287 ();
 fill_1 FILLER_87_301 ();
 fill_2 FILLER_87_327 ();
 fill_2 FILLER_87_346 ();
 fill_1 FILLER_87_348 ();
 fill_1 FILLER_87_365 ();
 fill_2 FILLER_87_390 ();
 fill_2 FILLER_87_399 ();
 fill_2 FILLER_87_408 ();
 fill_2 FILLER_87_419 ();
 fill_4 FILLER_87_429 ();
 fill_1 FILLER_87_444 ();
 fill_2 FILLER_87_479 ();
 fill_1 FILLER_87_576 ();
 fill_1 FILLER_87_597 ();
 fill_4 FILLER_87_629 ();
 fill_1 FILLER_87_633 ();
 fill_1 FILLER_87_659 ();
 fill_1 FILLER_87_671 ();
 fill_2 FILLER_87_682 ();
 fill_2 FILLER_87_696 ();
 fill_1 FILLER_87_698 ();
 fill_2 FILLER_87_719 ();
 fill_1 FILLER_87_721 ();
 fill_2 FILLER_87_725 ();
 fill_1 FILLER_87_727 ();
 fill_4 FILLER_87_733 ();
 fill_4 FILLER_87_759 ();
 fill_2 FILLER_87_763 ();
 fill_1 FILLER_87_765 ();
 fill_4 FILLER_87_777 ();
 fill_2 FILLER_87_781 ();
 fill_1 FILLER_87_783 ();
 decap_12 FILLER_87_841 ();
 decap_12 FILLER_87_853 ();
 decap_12 FILLER_87_865 ();
 decap_12 FILLER_87_877 ();
 fill_4 FILLER_87_889 ();
 fill_2 FILLER_87_893 ();
 fill_1 FILLER_87_895 ();
 decap_12 FILLER_87_897 ();
 decap_12 FILLER_87_909 ();
 decap_12 FILLER_87_921 ();
 decap_12 FILLER_87_933 ();
 fill_4 FILLER_87_945 ();
 fill_2 FILLER_87_949 ();
 fill_1 FILLER_87_951 ();
 decap_12 FILLER_87_953 ();
 decap_12 FILLER_87_965 ();
 decap_12 FILLER_87_977 ();
 decap_12 FILLER_87_989 ();
 fill_4 FILLER_87_1001 ();
 fill_2 FILLER_87_1005 ();
 fill_1 FILLER_87_1007 ();
 decap_12 FILLER_87_1009 ();
 decap_12 FILLER_87_1021 ();
 fill_4 FILLER_87_1033 ();
 fill_1 FILLER_87_1037 ();
 fill_4 FILLER_88_3 ();
 fill_1 FILLER_88_7 ();
 fill_2 FILLER_88_15 ();
 fill_1 FILLER_88_17 ();
 fill_4 FILLER_88_59 ();
 fill_2 FILLER_88_63 ();
 fill_8 FILLER_88_74 ();
 fill_2 FILLER_88_82 ();
 fill_2 FILLER_88_92 ();
 fill_1 FILLER_88_132 ();
 fill_4 FILLER_88_150 ();
 fill_8 FILLER_88_161 ();
 fill_2 FILLER_88_169 ();
 fill_2 FILLER_88_194 ();
 fill_1 FILLER_88_197 ();
 fill_1 FILLER_88_205 ();
 fill_1 FILLER_88_238 ();
 fill_2 FILLER_88_249 ();
 fill_1 FILLER_88_251 ();
 fill_2 FILLER_88_259 ();
 fill_1 FILLER_88_273 ();
 fill_4 FILLER_88_304 ();
 fill_4 FILLER_88_309 ();
 fill_1 FILLER_88_313 ();
 fill_4 FILLER_88_323 ();
 fill_1 FILLER_88_334 ();
 fill_2 FILLER_88_344 ();
 fill_1 FILLER_88_346 ();
 fill_1 FILLER_88_363 ();
 fill_2 FILLER_88_372 ();
 fill_2 FILLER_88_381 ();
 fill_1 FILLER_88_383 ();
 fill_1 FILLER_88_393 ();
 fill_2 FILLER_88_404 ();
 fill_1 FILLER_88_406 ();
 fill_4 FILLER_88_413 ();
 fill_2 FILLER_88_417 ();
 fill_1 FILLER_88_419 ();
 fill_4 FILLER_88_421 ();
 fill_4 FILLER_88_431 ();
 fill_2 FILLER_88_435 ();
 fill_1 FILLER_88_437 ();
 fill_2 FILLER_88_448 ();
 fill_1 FILLER_88_450 ();
 fill_1 FILLER_88_457 ();
 fill_2 FILLER_88_474 ();
 fill_2 FILLER_88_477 ();
 fill_1 FILLER_88_486 ();
 fill_1 FILLER_88_509 ();
 fill_2 FILLER_88_530 ();
 fill_4 FILLER_88_539 ();
 fill_2 FILLER_88_561 ();
 fill_1 FILLER_88_563 ();
 fill_2 FILLER_88_569 ();
 fill_4 FILLER_88_581 ();
 fill_8 FILLER_88_589 ();
 fill_2 FILLER_88_602 ();
 fill_1 FILLER_88_609 ();
 fill_2 FILLER_88_618 ();
 fill_1 FILLER_88_620 ();
 fill_4 FILLER_88_627 ();
 fill_1 FILLER_88_631 ();
 fill_4 FILLER_88_639 ();
 fill_1 FILLER_88_643 ();
 fill_8 FILLER_88_645 ();
 fill_8 FILLER_88_662 ();
 fill_2 FILLER_88_670 ();
 fill_1 FILLER_88_672 ();
 fill_4 FILLER_88_730 ();
 fill_1 FILLER_88_734 ();
 fill_4 FILLER_88_757 ();
 fill_1 FILLER_88_761 ();
 fill_2 FILLER_88_782 ();
 fill_1 FILLER_88_784 ();
 fill_2 FILLER_88_801 ();
 fill_1 FILLER_88_803 ();
 fill_4 FILLER_88_813 ();
 fill_2 FILLER_88_817 ();
 decap_12 FILLER_88_848 ();
 fill_8 FILLER_88_860 ();
 decap_12 FILLER_88_869 ();
 decap_12 FILLER_88_881 ();
 decap_12 FILLER_88_893 ();
 decap_12 FILLER_88_905 ();
 fill_4 FILLER_88_917 ();
 fill_2 FILLER_88_921 ();
 fill_1 FILLER_88_923 ();
 decap_12 FILLER_88_925 ();
 decap_12 FILLER_88_937 ();
 decap_12 FILLER_88_949 ();
 decap_12 FILLER_88_961 ();
 fill_4 FILLER_88_973 ();
 fill_2 FILLER_88_977 ();
 fill_1 FILLER_88_979 ();
 decap_12 FILLER_88_981 ();
 decap_12 FILLER_88_993 ();
 decap_12 FILLER_88_1005 ();
 decap_12 FILLER_88_1017 ();
 fill_4 FILLER_88_1029 ();
 fill_2 FILLER_88_1033 ();
 fill_1 FILLER_88_1035 ();
 fill_1 FILLER_88_1037 ();
 fill_1 FILLER_89_27 ();
 fill_4 FILLER_89_50 ();
 fill_2 FILLER_89_54 ();
 fill_1 FILLER_89_75 ();
 fill_1 FILLER_89_95 ();
 fill_1 FILLER_89_113 ();
 fill_4 FILLER_89_146 ();
 fill_1 FILLER_89_150 ();
 fill_1 FILLER_89_167 ();
 fill_1 FILLER_89_169 ();
 fill_4 FILLER_89_195 ();
 fill_1 FILLER_89_199 ();
 fill_2 FILLER_89_215 ();
 fill_4 FILLER_89_232 ();
 fill_2 FILLER_89_236 ();
 fill_1 FILLER_89_288 ();
 fill_2 FILLER_89_302 ();
 fill_8 FILLER_89_337 ();
 fill_4 FILLER_89_361 ();
 fill_1 FILLER_89_365 ();
 fill_2 FILLER_89_389 ();
 fill_1 FILLER_89_391 ();
 fill_4 FILLER_89_393 ();
 fill_2 FILLER_89_404 ();
 fill_2 FILLER_89_416 ();
 fill_1 FILLER_89_437 ();
 fill_1 FILLER_89_447 ();
 fill_2 FILLER_89_453 ();
 fill_2 FILLER_89_465 ();
 fill_2 FILLER_89_482 ();
 fill_1 FILLER_89_513 ();
 fill_2 FILLER_89_558 ();
 fill_1 FILLER_89_561 ();
 fill_4 FILLER_89_574 ();
 fill_2 FILLER_89_578 ();
 fill_8 FILLER_89_587 ();
 fill_1 FILLER_89_595 ();
 fill_1 FILLER_89_615 ();
 fill_8 FILLER_89_634 ();
 fill_4 FILLER_89_646 ();
 fill_2 FILLER_89_650 ();
 fill_1 FILLER_89_652 ();
 fill_2 FILLER_89_657 ();
 fill_1 FILLER_89_680 ();
 fill_4 FILLER_89_684 ();
 fill_1 FILLER_89_688 ();
 fill_4 FILLER_89_699 ();
 fill_1 FILLER_89_703 ();
 fill_2 FILLER_89_726 ();
 fill_4 FILLER_89_777 ();
 fill_2 FILLER_89_781 ();
 fill_1 FILLER_89_783 ();
 fill_4 FILLER_89_794 ();
 fill_2 FILLER_89_798 ();
 decap_12 FILLER_89_857 ();
 decap_12 FILLER_89_869 ();
 decap_12 FILLER_89_881 ();
 fill_2 FILLER_89_893 ();
 fill_1 FILLER_89_895 ();
 decap_12 FILLER_89_897 ();
 decap_12 FILLER_89_909 ();
 decap_12 FILLER_89_921 ();
 decap_12 FILLER_89_933 ();
 fill_4 FILLER_89_945 ();
 fill_2 FILLER_89_949 ();
 fill_1 FILLER_89_951 ();
 decap_12 FILLER_89_953 ();
 decap_12 FILLER_89_965 ();
 decap_12 FILLER_89_977 ();
 decap_12 FILLER_89_989 ();
 fill_4 FILLER_89_1001 ();
 fill_2 FILLER_89_1005 ();
 fill_1 FILLER_89_1007 ();
 decap_12 FILLER_89_1009 ();
 decap_12 FILLER_89_1021 ();
 fill_4 FILLER_89_1033 ();
 fill_1 FILLER_89_1037 ();
 fill_4 FILLER_90_3 ();
 fill_2 FILLER_90_7 ();
 fill_1 FILLER_90_9 ();
 decap_12 FILLER_90_29 ();
 fill_1 FILLER_90_41 ();
 fill_4 FILLER_90_51 ();
 fill_2 FILLER_90_55 ();
 fill_2 FILLER_90_64 ();
 fill_1 FILLER_90_66 ();
 fill_4 FILLER_90_71 ();
 fill_2 FILLER_90_75 ();
 fill_2 FILLER_90_81 ();
 fill_1 FILLER_90_83 ();
 fill_8 FILLER_90_89 ();
 fill_4 FILLER_90_113 ();
 fill_2 FILLER_90_117 ();
 decap_12 FILLER_90_126 ();
 fill_2 FILLER_90_138 ();
 fill_2 FILLER_90_157 ();
 fill_1 FILLER_90_159 ();
 fill_4 FILLER_90_169 ();
 fill_1 FILLER_90_173 ();
 fill_2 FILLER_90_188 ();
 fill_2 FILLER_90_209 ();
 fill_2 FILLER_90_220 ();
 fill_4 FILLER_90_235 ();
 fill_2 FILLER_90_246 ();
 fill_8 FILLER_90_260 ();
 fill_1 FILLER_90_287 ();
 fill_4 FILLER_90_318 ();
 fill_1 FILLER_90_329 ();
 decap_12 FILLER_90_335 ();
 fill_2 FILLER_90_347 ();
 fill_4 FILLER_90_358 ();
 fill_2 FILLER_90_362 ();
 fill_2 FILLER_90_372 ();
 fill_2 FILLER_90_399 ();
 fill_1 FILLER_90_401 ();
 fill_2 FILLER_90_410 ();
 fill_1 FILLER_90_412 ();
 fill_1 FILLER_90_421 ();
 fill_2 FILLER_90_429 ();
 fill_2 FILLER_90_438 ();
 fill_1 FILLER_90_440 ();
 fill_1 FILLER_90_468 ();
 fill_1 FILLER_90_497 ();
 fill_1 FILLER_90_504 ();
 fill_1 FILLER_90_513 ();
 fill_2 FILLER_90_529 ();
 fill_1 FILLER_90_531 ();
 fill_4 FILLER_90_558 ();
 fill_1 FILLER_90_562 ();
 decap_12 FILLER_90_572 ();
 fill_4 FILLER_90_584 ();
 fill_2 FILLER_90_600 ();
 decap_12 FILLER_90_608 ();
 fill_2 FILLER_90_620 ();
 fill_1 FILLER_90_643 ();
 fill_2 FILLER_90_656 ();
 fill_1 FILLER_90_658 ();
 fill_2 FILLER_90_672 ();
 fill_2 FILLER_90_681 ();
 fill_4 FILLER_90_722 ();
 fill_2 FILLER_90_726 ();
 fill_2 FILLER_90_737 ();
 fill_1 FILLER_90_739 ();
 fill_4 FILLER_90_806 ();
 fill_2 FILLER_90_810 ();
 decap_12 FILLER_90_846 ();
 fill_8 FILLER_90_858 ();
 fill_2 FILLER_90_866 ();
 decap_12 FILLER_90_869 ();
 decap_12 FILLER_90_881 ();
 decap_12 FILLER_90_893 ();
 decap_12 FILLER_90_905 ();
 fill_4 FILLER_90_917 ();
 fill_2 FILLER_90_921 ();
 fill_1 FILLER_90_923 ();
 decap_12 FILLER_90_925 ();
 decap_12 FILLER_90_937 ();
 decap_12 FILLER_90_949 ();
 decap_12 FILLER_90_961 ();
 fill_4 FILLER_90_973 ();
 fill_2 FILLER_90_977 ();
 fill_1 FILLER_90_979 ();
 decap_12 FILLER_90_981 ();
 decap_12 FILLER_90_993 ();
 decap_12 FILLER_90_1005 ();
 decap_12 FILLER_90_1017 ();
 fill_4 FILLER_90_1029 ();
 fill_1 FILLER_90_1037 ();
 fill_1 FILLER_91_3 ();
 fill_2 FILLER_91_21 ();
 fill_2 FILLER_91_36 ();
 fill_2 FILLER_91_53 ();
 fill_1 FILLER_91_55 ();
 fill_4 FILLER_91_65 ();
 fill_2 FILLER_91_69 ();
 fill_1 FILLER_91_71 ();
 fill_2 FILLER_91_83 ();
 fill_1 FILLER_91_85 ();
 fill_1 FILLER_91_111 ();
 fill_1 FILLER_91_113 ();
 fill_8 FILLER_91_135 ();
 fill_4 FILLER_91_164 ();
 fill_4 FILLER_91_202 ();
 fill_8 FILLER_91_214 ();
 fill_2 FILLER_91_222 ();
 fill_2 FILLER_91_225 ();
 fill_4 FILLER_91_231 ();
 fill_1 FILLER_91_235 ();
 fill_2 FILLER_91_281 ();
 fill_1 FILLER_91_283 ();
 fill_2 FILLER_91_316 ();
 fill_2 FILLER_91_334 ();
 fill_1 FILLER_91_337 ();
 fill_1 FILLER_91_354 ();
 fill_2 FILLER_91_393 ();
 fill_1 FILLER_91_395 ();
 fill_4 FILLER_91_399 ();
 fill_2 FILLER_91_403 ();
 fill_4 FILLER_91_421 ();
 fill_1 FILLER_91_428 ();
 fill_2 FILLER_91_432 ();
 fill_1 FILLER_91_434 ();
 fill_4 FILLER_91_438 ();
 fill_2 FILLER_91_476 ();
 fill_1 FILLER_91_492 ();
 fill_2 FILLER_91_501 ();
 fill_1 FILLER_91_503 ();
 fill_1 FILLER_91_533 ();
 fill_2 FILLER_91_575 ();
 fill_1 FILLER_91_577 ();
 fill_2 FILLER_91_587 ();
 fill_4 FILLER_91_595 ();
 fill_1 FILLER_91_599 ();
 fill_8 FILLER_91_606 ();
 fill_2 FILLER_91_614 ();
 decap_12 FILLER_91_624 ();
 decap_12 FILLER_91_636 ();
 fill_2 FILLER_91_662 ();
 fill_4 FILLER_91_673 ();
 fill_2 FILLER_91_677 ();
 fill_1 FILLER_91_688 ();
 fill_4 FILLER_91_697 ();
 fill_2 FILLER_91_701 ();
 fill_4 FILLER_91_708 ();
 fill_2 FILLER_91_781 ();
 fill_1 FILLER_91_783 ();
 fill_4 FILLER_91_785 ();
 fill_2 FILLER_91_789 ();
 fill_1 FILLER_91_808 ();
 fill_4 FILLER_91_827 ();
 decap_12 FILLER_91_841 ();
 decap_12 FILLER_91_853 ();
 decap_12 FILLER_91_865 ();
 decap_12 FILLER_91_877 ();
 fill_4 FILLER_91_889 ();
 fill_2 FILLER_91_893 ();
 fill_1 FILLER_91_895 ();
 decap_12 FILLER_91_897 ();
 decap_12 FILLER_91_909 ();
 decap_12 FILLER_91_921 ();
 decap_12 FILLER_91_933 ();
 fill_4 FILLER_91_945 ();
 fill_2 FILLER_91_949 ();
 fill_1 FILLER_91_951 ();
 decap_12 FILLER_91_953 ();
 decap_12 FILLER_91_965 ();
 decap_12 FILLER_91_977 ();
 decap_12 FILLER_91_989 ();
 fill_4 FILLER_91_1001 ();
 fill_2 FILLER_91_1005 ();
 fill_1 FILLER_91_1007 ();
 decap_12 FILLER_91_1009 ();
 decap_12 FILLER_91_1021 ();
 fill_4 FILLER_91_1033 ();
 fill_1 FILLER_91_1037 ();
 fill_4 FILLER_92_3 ();
 fill_2 FILLER_92_7 ();
 fill_4 FILLER_92_24 ();
 fill_4 FILLER_92_41 ();
 fill_2 FILLER_92_45 ();
 fill_2 FILLER_92_55 ();
 fill_1 FILLER_92_57 ();
 fill_2 FILLER_92_81 ();
 fill_1 FILLER_92_83 ();
 fill_1 FILLER_92_104 ();
 fill_8 FILLER_92_121 ();
 fill_1 FILLER_92_129 ();
 fill_1 FILLER_92_139 ();
 fill_4 FILLER_92_150 ();
 fill_4 FILLER_92_163 ();
 fill_2 FILLER_92_172 ();
 fill_2 FILLER_92_187 ();
 fill_1 FILLER_92_189 ();
 fill_1 FILLER_92_197 ();
 fill_4 FILLER_92_212 ();
 fill_1 FILLER_92_216 ();
 fill_1 FILLER_92_224 ();
 fill_2 FILLER_92_299 ();
 fill_2 FILLER_92_318 ();
 fill_1 FILLER_92_372 ();
 decap_12 FILLER_92_389 ();
 fill_2 FILLER_92_417 ();
 fill_1 FILLER_92_419 ();
 fill_2 FILLER_92_429 ();
 fill_1 FILLER_92_497 ();
 fill_1 FILLER_92_546 ();
 fill_2 FILLER_92_558 ();
 fill_2 FILLER_92_567 ();
 fill_1 FILLER_92_569 ();
 fill_4 FILLER_92_577 ();
 fill_1 FILLER_92_596 ();
 fill_2 FILLER_92_609 ();
 fill_1 FILLER_92_611 ();
 fill_2 FILLER_92_626 ();
 fill_4 FILLER_92_637 ();
 fill_2 FILLER_92_641 ();
 fill_1 FILLER_92_643 ();
 fill_1 FILLER_92_652 ();
 fill_2 FILLER_92_658 ();
 fill_1 FILLER_92_667 ();
 fill_2 FILLER_92_683 ();
 fill_2 FILLER_92_698 ();
 fill_2 FILLER_92_717 ();
 fill_1 FILLER_92_728 ();
 fill_4 FILLER_92_736 ();
 fill_4 FILLER_92_757 ();
 fill_1 FILLER_92_761 ();
 fill_1 FILLER_92_778 ();
 fill_1 FILLER_92_811 ();
 decap_12 FILLER_92_845 ();
 fill_8 FILLER_92_857 ();
 fill_2 FILLER_92_865 ();
 fill_1 FILLER_92_867 ();
 decap_12 FILLER_92_869 ();
 decap_12 FILLER_92_881 ();
 decap_12 FILLER_92_893 ();
 decap_12 FILLER_92_905 ();
 fill_4 FILLER_92_917 ();
 fill_2 FILLER_92_921 ();
 fill_1 FILLER_92_923 ();
 decap_12 FILLER_92_925 ();
 decap_12 FILLER_92_937 ();
 decap_12 FILLER_92_949 ();
 decap_12 FILLER_92_961 ();
 fill_4 FILLER_92_973 ();
 fill_2 FILLER_92_977 ();
 fill_1 FILLER_92_979 ();
 decap_12 FILLER_92_981 ();
 decap_12 FILLER_92_993 ();
 decap_12 FILLER_92_1005 ();
 decap_12 FILLER_92_1017 ();
 fill_4 FILLER_92_1029 ();
 fill_2 FILLER_92_1033 ();
 fill_1 FILLER_92_1035 ();
 fill_1 FILLER_92_1037 ();
 fill_1 FILLER_93_22 ();
 fill_1 FILLER_93_47 ();
 fill_1 FILLER_93_57 ();
 fill_2 FILLER_93_83 ();
 fill_2 FILLER_93_110 ();
 fill_2 FILLER_93_126 ();
 fill_1 FILLER_93_144 ();
 fill_2 FILLER_93_213 ();
 fill_1 FILLER_93_215 ();
 fill_2 FILLER_93_222 ();
 fill_2 FILLER_93_231 ();
 fill_1 FILLER_93_263 ();
 fill_2 FILLER_93_271 ();
 fill_2 FILLER_93_281 ();
 fill_1 FILLER_93_283 ();
 fill_1 FILLER_93_353 ();
 fill_4 FILLER_93_363 ();
 fill_2 FILLER_93_390 ();
 fill_8 FILLER_93_431 ();
 fill_1 FILLER_93_444 ();
 fill_2 FILLER_93_449 ();
 fill_1 FILLER_93_470 ();
 fill_1 FILLER_93_479 ();
 fill_2 FILLER_93_489 ();
 fill_2 FILLER_93_498 ();
 fill_4 FILLER_93_542 ();
 fill_2 FILLER_93_561 ();
 decap_12 FILLER_93_571 ();
 decap_12 FILLER_93_583 ();
 fill_1 FILLER_93_595 ();
 fill_1 FILLER_93_601 ();
 fill_4 FILLER_93_610 ();
 fill_2 FILLER_93_614 ();
 fill_2 FILLER_93_623 ();
 fill_1 FILLER_93_625 ();
 fill_2 FILLER_93_629 ();
 fill_1 FILLER_93_631 ();
 fill_4 FILLER_93_680 ();
 fill_2 FILLER_93_684 ();
 fill_4 FILLER_93_701 ();
 fill_2 FILLER_93_705 ();
 fill_1 FILLER_93_716 ();
 fill_2 FILLER_93_726 ();
 fill_1 FILLER_93_729 ();
 fill_1 FILLER_93_747 ();
 fill_2 FILLER_93_766 ();
 fill_1 FILLER_93_777 ();
 fill_2 FILLER_93_794 ();
 fill_2 FILLER_93_805 ();
 fill_1 FILLER_93_824 ();
 fill_2 FILLER_93_837 ();
 fill_1 FILLER_93_839 ();
 decap_12 FILLER_93_841 ();
 decap_12 FILLER_93_853 ();
 decap_12 FILLER_93_865 ();
 decap_12 FILLER_93_877 ();
 fill_4 FILLER_93_889 ();
 fill_2 FILLER_93_893 ();
 fill_1 FILLER_93_895 ();
 decap_12 FILLER_93_897 ();
 decap_12 FILLER_93_909 ();
 decap_12 FILLER_93_921 ();
 decap_12 FILLER_93_933 ();
 fill_4 FILLER_93_945 ();
 fill_2 FILLER_93_949 ();
 fill_1 FILLER_93_951 ();
 decap_12 FILLER_93_953 ();
 decap_12 FILLER_93_965 ();
 decap_12 FILLER_93_977 ();
 decap_12 FILLER_93_989 ();
 fill_4 FILLER_93_1001 ();
 fill_2 FILLER_93_1005 ();
 fill_1 FILLER_93_1007 ();
 decap_12 FILLER_93_1009 ();
 decap_12 FILLER_93_1021 ();
 fill_4 FILLER_93_1033 ();
 fill_1 FILLER_93_1037 ();
 fill_4 FILLER_94_3 ();
 fill_2 FILLER_94_7 ();
 fill_4 FILLER_94_21 ();
 fill_2 FILLER_94_25 ();
 fill_1 FILLER_94_27 ();
 fill_4 FILLER_94_29 ();
 fill_1 FILLER_94_33 ();
 fill_1 FILLER_94_53 ();
 fill_1 FILLER_94_83 ();
 fill_4 FILLER_94_85 ();
 fill_2 FILLER_94_89 ();
 fill_1 FILLER_94_91 ();
 fill_4 FILLER_94_101 ();
 fill_2 FILLER_94_105 ();
 fill_2 FILLER_94_137 ();
 fill_1 FILLER_94_139 ();
 fill_2 FILLER_94_152 ();
 fill_1 FILLER_94_154 ();
 fill_4 FILLER_94_164 ();
 fill_2 FILLER_94_168 ();
 fill_4 FILLER_94_177 ();
 fill_2 FILLER_94_187 ();
 fill_1 FILLER_94_210 ();
 fill_1 FILLER_94_218 ();
 fill_2 FILLER_94_305 ();
 fill_1 FILLER_94_307 ();
 fill_1 FILLER_94_309 ();
 fill_2 FILLER_94_319 ();
 fill_1 FILLER_94_321 ();
 fill_2 FILLER_94_335 ();
 fill_1 FILLER_94_337 ();
 fill_1 FILLER_94_363 ();
 fill_2 FILLER_94_377 ();
 fill_4 FILLER_94_400 ();
 fill_4 FILLER_94_416 ();
 fill_4 FILLER_94_424 ();
 fill_2 FILLER_94_428 ();
 fill_1 FILLER_94_430 ();
 fill_1 FILLER_94_475 ();
 fill_2 FILLER_94_514 ();
 fill_1 FILLER_94_551 ();
 fill_2 FILLER_94_567 ();
 fill_2 FILLER_94_577 ();
 fill_2 FILLER_94_586 ();
 fill_8 FILLER_94_597 ();
 fill_1 FILLER_94_605 ();
 fill_4 FILLER_94_629 ();
 fill_1 FILLER_94_633 ();
 fill_4 FILLER_94_639 ();
 fill_1 FILLER_94_643 ();
 fill_4 FILLER_94_645 ();
 fill_2 FILLER_94_649 ();
 fill_1 FILLER_94_651 ();
 fill_2 FILLER_94_669 ();
 fill_1 FILLER_94_671 ();
 fill_2 FILLER_94_676 ();
 fill_1 FILLER_94_678 ();
 fill_4 FILLER_94_695 ();
 fill_1 FILLER_94_699 ();
 fill_4 FILLER_94_749 ();
 fill_1 FILLER_94_786 ();
 fill_2 FILLER_94_794 ();
 fill_1 FILLER_94_796 ();
 fill_2 FILLER_94_818 ();
 decap_12 FILLER_94_845 ();
 fill_8 FILLER_94_857 ();
 fill_2 FILLER_94_865 ();
 fill_1 FILLER_94_867 ();
 decap_12 FILLER_94_869 ();
 decap_12 FILLER_94_881 ();
 decap_12 FILLER_94_893 ();
 decap_12 FILLER_94_905 ();
 fill_4 FILLER_94_917 ();
 fill_2 FILLER_94_921 ();
 fill_1 FILLER_94_923 ();
 decap_12 FILLER_94_925 ();
 decap_12 FILLER_94_937 ();
 decap_12 FILLER_94_949 ();
 decap_12 FILLER_94_961 ();
 fill_4 FILLER_94_973 ();
 fill_2 FILLER_94_977 ();
 fill_1 FILLER_94_979 ();
 decap_12 FILLER_94_981 ();
 decap_12 FILLER_94_993 ();
 decap_12 FILLER_94_1005 ();
 decap_12 FILLER_94_1017 ();
 fill_4 FILLER_94_1029 ();
 fill_2 FILLER_94_1033 ();
 fill_1 FILLER_94_1035 ();
 fill_1 FILLER_94_1037 ();
 fill_2 FILLER_95_3 ();
 fill_1 FILLER_95_25 ();
 fill_1 FILLER_95_48 ();
 fill_4 FILLER_95_52 ();
 fill_2 FILLER_95_122 ();
 fill_2 FILLER_95_152 ();
 fill_2 FILLER_95_161 ();
 fill_1 FILLER_95_163 ();
 fill_4 FILLER_95_202 ();
 fill_1 FILLER_95_209 ();
 fill_2 FILLER_95_216 ();
 fill_1 FILLER_95_218 ();
 fill_1 FILLER_95_223 ();
 fill_2 FILLER_95_277 ();
 fill_1 FILLER_95_279 ();
 fill_2 FILLER_95_315 ();
 fill_1 FILLER_95_317 ();
 fill_4 FILLER_95_327 ();
 fill_1 FILLER_95_331 ();
 fill_1 FILLER_95_371 ();
 fill_4 FILLER_95_388 ();
 fill_4 FILLER_95_393 ();
 fill_1 FILLER_95_397 ();
 fill_2 FILLER_95_418 ();
 fill_1 FILLER_95_427 ();
 fill_2 FILLER_95_458 ();
 fill_1 FILLER_95_469 ();
 fill_2 FILLER_95_483 ();
 fill_1 FILLER_95_485 ();
 fill_4 FILLER_95_489 ();
 fill_1 FILLER_95_493 ();
 fill_2 FILLER_95_505 ();
 fill_1 FILLER_95_507 ();
 fill_1 FILLER_95_529 ();
 fill_2 FILLER_95_546 ();
 fill_1 FILLER_95_559 ();
 fill_8 FILLER_95_583 ();
 fill_2 FILLER_95_591 ();
 fill_1 FILLER_95_593 ();
 fill_4 FILLER_95_623 ();
 fill_2 FILLER_95_634 ();
 fill_2 FILLER_95_647 ();
 fill_1 FILLER_95_668 ();
 fill_4 FILLER_95_680 ();
 fill_1 FILLER_95_684 ();
 fill_2 FILLER_95_688 ();
 fill_4 FILLER_95_697 ();
 fill_1 FILLER_95_701 ();
 decap_12 FILLER_95_714 ();
 fill_2 FILLER_95_726 ();
 fill_4 FILLER_95_772 ();
 fill_2 FILLER_95_781 ();
 fill_1 FILLER_95_783 ();
 fill_1 FILLER_95_785 ();
 fill_2 FILLER_95_814 ();
 decap_12 FILLER_95_841 ();
 decap_12 FILLER_95_853 ();
 decap_12 FILLER_95_865 ();
 decap_12 FILLER_95_877 ();
 fill_4 FILLER_95_889 ();
 fill_2 FILLER_95_893 ();
 fill_1 FILLER_95_895 ();
 decap_12 FILLER_95_897 ();
 decap_12 FILLER_95_909 ();
 decap_12 FILLER_95_921 ();
 decap_12 FILLER_95_933 ();
 fill_4 FILLER_95_945 ();
 fill_2 FILLER_95_949 ();
 fill_1 FILLER_95_951 ();
 decap_12 FILLER_95_953 ();
 decap_12 FILLER_95_965 ();
 decap_12 FILLER_95_977 ();
 decap_12 FILLER_95_989 ();
 fill_4 FILLER_95_1001 ();
 fill_2 FILLER_95_1005 ();
 fill_1 FILLER_95_1007 ();
 decap_12 FILLER_95_1009 ();
 decap_12 FILLER_95_1021 ();
 fill_4 FILLER_95_1033 ();
 fill_1 FILLER_95_1037 ();
 fill_2 FILLER_96_3 ();
 fill_2 FILLER_96_72 ();
 fill_1 FILLER_96_74 ();
 fill_2 FILLER_96_85 ();
 fill_1 FILLER_96_101 ();
 fill_2 FILLER_96_141 ();
 fill_1 FILLER_96_143 ();
 fill_2 FILLER_96_170 ();
 fill_1 FILLER_96_172 ();
 fill_1 FILLER_96_197 ();
 fill_2 FILLER_96_206 ();
 fill_2 FILLER_96_236 ();
 fill_1 FILLER_96_238 ();
 fill_1 FILLER_96_251 ();
 fill_2 FILLER_96_267 ();
 fill_1 FILLER_96_269 ();
 fill_1 FILLER_96_300 ();
 fill_1 FILLER_96_309 ();
 fill_1 FILLER_96_330 ();
 fill_1 FILLER_96_347 ();
 fill_1 FILLER_96_365 ();
 fill_2 FILLER_96_418 ();
 fill_1 FILLER_96_428 ();
 fill_1 FILLER_96_438 ();
 fill_1 FILLER_96_442 ();
 fill_2 FILLER_96_450 ();
 fill_1 FILLER_96_468 ();
 fill_1 FILLER_96_477 ();
 fill_4 FILLER_96_498 ();
 fill_1 FILLER_96_502 ();
 fill_2 FILLER_96_510 ();
 fill_1 FILLER_96_512 ();
 fill_2 FILLER_96_520 ();
 fill_4 FILLER_96_527 ();
 fill_1 FILLER_96_531 ();
 fill_1 FILLER_96_533 ();
 fill_1 FILLER_96_546 ();
 fill_1 FILLER_96_574 ();
 fill_2 FILLER_96_586 ();
 decap_12 FILLER_96_589 ();
 decap_12 FILLER_96_604 ();
 fill_4 FILLER_96_616 ();
 fill_1 FILLER_96_620 ();
 fill_1 FILLER_96_627 ();
 fill_4 FILLER_96_640 ();
 fill_4 FILLER_96_652 ();
 fill_1 FILLER_96_664 ();
 fill_1 FILLER_96_674 ();
 fill_1 FILLER_96_679 ();
 fill_2 FILLER_96_698 ();
 fill_8 FILLER_96_736 ();
 fill_2 FILLER_96_753 ();
 fill_1 FILLER_96_755 ();
 fill_8 FILLER_96_765 ();
 fill_1 FILLER_96_781 ();
 fill_1 FILLER_96_804 ();
 fill_4 FILLER_96_813 ();
 fill_2 FILLER_96_827 ();
 decap_12 FILLER_96_838 ();
 decap_12 FILLER_96_850 ();
 fill_4 FILLER_96_862 ();
 fill_2 FILLER_96_866 ();
 decap_12 FILLER_96_869 ();
 decap_12 FILLER_96_881 ();
 decap_12 FILLER_96_893 ();
 decap_12 FILLER_96_905 ();
 fill_4 FILLER_96_917 ();
 fill_2 FILLER_96_921 ();
 fill_1 FILLER_96_923 ();
 decap_12 FILLER_96_925 ();
 decap_12 FILLER_96_937 ();
 decap_12 FILLER_96_949 ();
 decap_12 FILLER_96_961 ();
 fill_4 FILLER_96_973 ();
 fill_2 FILLER_96_977 ();
 fill_1 FILLER_96_979 ();
 decap_12 FILLER_96_981 ();
 decap_12 FILLER_96_993 ();
 decap_12 FILLER_96_1005 ();
 decap_12 FILLER_96_1017 ();
 fill_4 FILLER_96_1029 ();
 fill_2 FILLER_96_1033 ();
 fill_1 FILLER_96_1035 ();
 fill_1 FILLER_96_1037 ();
 fill_2 FILLER_97_3 ();
 fill_4 FILLER_97_14 ();
 fill_1 FILLER_97_18 ();
 fill_4 FILLER_97_31 ();
 fill_2 FILLER_97_35 ();
 fill_2 FILLER_97_53 ();
 fill_1 FILLER_97_55 ();
 fill_2 FILLER_97_110 ();
 fill_1 FILLER_97_129 ();
 fill_2 FILLER_97_155 ();
 fill_4 FILLER_97_164 ();
 fill_1 FILLER_97_169 ();
 fill_2 FILLER_97_183 ();
 fill_1 FILLER_97_219 ();
 fill_1 FILLER_97_260 ();
 fill_1 FILLER_97_279 ();
 fill_4 FILLER_97_281 ();
 fill_2 FILLER_97_285 ();
 fill_1 FILLER_97_287 ();
 fill_1 FILLER_97_294 ();
 fill_1 FILLER_97_317 ();
 fill_2 FILLER_97_327 ();
 fill_2 FILLER_97_357 ();
 fill_4 FILLER_97_375 ();
 fill_4 FILLER_97_388 ();
 fill_8 FILLER_97_393 ();
 fill_1 FILLER_97_447 ();
 fill_2 FILLER_97_472 ();
 fill_4 FILLER_97_482 ();
 fill_1 FILLER_97_486 ();
 fill_2 FILLER_97_501 ();
 fill_1 FILLER_97_503 ();
 fill_4 FILLER_97_543 ();
 fill_2 FILLER_97_547 ();
 fill_4 FILLER_97_561 ();
 fill_2 FILLER_97_565 ();
 fill_2 FILLER_97_575 ();
 fill_2 FILLER_97_584 ();
 fill_1 FILLER_97_605 ();
 fill_1 FILLER_97_609 ();
 fill_2 FILLER_97_613 ();
 fill_1 FILLER_97_615 ();
 fill_1 FILLER_97_617 ();
 fill_2 FILLER_97_624 ();
 fill_1 FILLER_97_626 ();
 fill_4 FILLER_97_631 ();
 fill_2 FILLER_97_635 ();
 fill_8 FILLER_97_643 ();
 fill_8 FILLER_97_663 ();
 fill_1 FILLER_97_671 ();
 fill_1 FILLER_97_689 ();
 fill_8 FILLER_97_698 ();
 fill_2 FILLER_97_706 ();
 fill_4 FILLER_97_723 ();
 fill_1 FILLER_97_727 ();
 fill_2 FILLER_97_729 ();
 fill_4 FILLER_97_773 ();
 fill_2 FILLER_97_777 ();
 fill_4 FILLER_97_785 ();
 fill_1 FILLER_97_789 ();
 fill_1 FILLER_97_806 ();
 fill_1 FILLER_97_822 ();
 fill_2 FILLER_97_838 ();
 decap_12 FILLER_97_846 ();
 decap_12 FILLER_97_858 ();
 decap_12 FILLER_97_870 ();
 decap_12 FILLER_97_882 ();
 fill_2 FILLER_97_894 ();
 decap_12 FILLER_97_897 ();
 decap_12 FILLER_97_909 ();
 decap_12 FILLER_97_921 ();
 decap_12 FILLER_97_933 ();
 fill_4 FILLER_97_945 ();
 fill_2 FILLER_97_949 ();
 fill_1 FILLER_97_951 ();
 decap_12 FILLER_97_953 ();
 decap_12 FILLER_97_965 ();
 decap_12 FILLER_97_977 ();
 decap_12 FILLER_97_989 ();
 fill_4 FILLER_97_1001 ();
 fill_2 FILLER_97_1005 ();
 fill_1 FILLER_97_1007 ();
 decap_12 FILLER_97_1009 ();
 decap_12 FILLER_97_1021 ();
 fill_4 FILLER_97_1033 ();
 fill_1 FILLER_97_1037 ();
 fill_2 FILLER_98_26 ();
 fill_1 FILLER_98_29 ();
 fill_4 FILLER_98_39 ();
 fill_2 FILLER_98_43 ();
 fill_4 FILLER_98_61 ();
 fill_1 FILLER_98_69 ();
 fill_4 FILLER_98_79 ();
 fill_1 FILLER_98_83 ();
 fill_2 FILLER_98_94 ();
 fill_4 FILLER_98_121 ();
 fill_2 FILLER_98_125 ();
 fill_4 FILLER_98_134 ();
 fill_2 FILLER_98_138 ();
 fill_1 FILLER_98_150 ();
 fill_1 FILLER_98_197 ();
 fill_1 FILLER_98_219 ();
 fill_1 FILLER_98_238 ();
 fill_4 FILLER_98_247 ();
 fill_1 FILLER_98_251 ();
 fill_1 FILLER_98_289 ();
 fill_2 FILLER_98_306 ();
 fill_4 FILLER_98_309 ();
 fill_2 FILLER_98_322 ();
 fill_2 FILLER_98_327 ();
 fill_1 FILLER_98_329 ();
 fill_4 FILLER_98_339 ();
 fill_2 FILLER_98_343 ();
 fill_1 FILLER_98_363 ();
 fill_4 FILLER_98_365 ();
 fill_2 FILLER_98_406 ();
 fill_2 FILLER_98_421 ();
 fill_4 FILLER_98_435 ();
 fill_2 FILLER_98_439 ();
 fill_8 FILLER_98_444 ();
 fill_2 FILLER_98_452 ();
 fill_4 FILLER_98_472 ();
 fill_8 FILLER_98_484 ();
 fill_1 FILLER_98_492 ();
 fill_1 FILLER_98_501 ();
 fill_2 FILLER_98_530 ();
 fill_4 FILLER_98_561 ();
 fill_1 FILLER_98_587 ();
 fill_1 FILLER_98_599 ();
 fill_1 FILLER_98_609 ();
 fill_2 FILLER_98_642 ();
 fill_2 FILLER_98_649 ();
 fill_4 FILLER_98_666 ();
 fill_1 FILLER_98_675 ();
 fill_1 FILLER_98_683 ();
 fill_2 FILLER_98_697 ();
 fill_1 FILLER_98_699 ();
 decap_12 FILLER_98_722 ();
 fill_4 FILLER_98_750 ();
 fill_2 FILLER_98_754 ();
 fill_4 FILLER_98_757 ();
 fill_1 FILLER_98_761 ();
 fill_2 FILLER_98_771 ();
 fill_4 FILLER_98_795 ();
 fill_1 FILLER_98_799 ();
 fill_8 FILLER_98_804 ();
 fill_2 FILLER_98_813 ();
 fill_1 FILLER_98_825 ();
 decap_12 FILLER_98_849 ();
 fill_4 FILLER_98_861 ();
 fill_2 FILLER_98_865 ();
 fill_1 FILLER_98_867 ();
 decap_12 FILLER_98_869 ();
 decap_12 FILLER_98_881 ();
 decap_12 FILLER_98_893 ();
 decap_12 FILLER_98_905 ();
 fill_4 FILLER_98_917 ();
 fill_2 FILLER_98_921 ();
 fill_1 FILLER_98_923 ();
 decap_12 FILLER_98_925 ();
 decap_12 FILLER_98_937 ();
 decap_12 FILLER_98_949 ();
 decap_12 FILLER_98_961 ();
 fill_4 FILLER_98_973 ();
 fill_2 FILLER_98_977 ();
 fill_1 FILLER_98_979 ();
 decap_12 FILLER_98_981 ();
 decap_12 FILLER_98_993 ();
 decap_12 FILLER_98_1005 ();
 decap_12 FILLER_98_1017 ();
 fill_4 FILLER_98_1029 ();
 fill_2 FILLER_98_1033 ();
 fill_1 FILLER_98_1035 ();
 fill_1 FILLER_98_1037 ();
 fill_4 FILLER_99_3 ();
 fill_1 FILLER_99_7 ();
 fill_1 FILLER_99_21 ();
 fill_2 FILLER_99_54 ();
 fill_2 FILLER_99_57 ();
 fill_1 FILLER_99_59 ();
 fill_4 FILLER_99_88 ();
 fill_1 FILLER_99_92 ();
 fill_2 FILLER_99_102 ();
 fill_1 FILLER_99_111 ();
 fill_1 FILLER_99_113 ();
 fill_2 FILLER_99_146 ();
 fill_2 FILLER_99_154 ();
 fill_1 FILLER_99_156 ();
 fill_4 FILLER_99_163 ();
 fill_1 FILLER_99_167 ();
 fill_8 FILLER_99_169 ();
 fill_1 FILLER_99_177 ();
 fill_2 FILLER_99_202 ();
 fill_2 FILLER_99_236 ();
 fill_1 FILLER_99_253 ();
 fill_2 FILLER_99_272 ();
 fill_1 FILLER_99_291 ();
 fill_4 FILLER_99_353 ();
 fill_2 FILLER_99_371 ();
 fill_2 FILLER_99_389 ();
 fill_1 FILLER_99_391 ();
 fill_2 FILLER_99_393 ();
 fill_1 FILLER_99_482 ();
 fill_1 FILLER_99_503 ();
 fill_4 FILLER_99_529 ();
 fill_2 FILLER_99_533 ();
 fill_1 FILLER_99_535 ();
 fill_2 FILLER_99_558 ();
 decap_12 FILLER_99_596 ();
 fill_8 FILLER_99_608 ();
 decap_12 FILLER_99_626 ();
 decap_12 FILLER_99_638 ();
 fill_8 FILLER_99_650 ();
 fill_4 FILLER_99_667 ();
 fill_1 FILLER_99_671 ();
 fill_2 FILLER_99_682 ();
 fill_1 FILLER_99_700 ();
 fill_4 FILLER_99_722 ();
 fill_2 FILLER_99_726 ();
 fill_8 FILLER_99_729 ();
 fill_2 FILLER_99_737 ();
 fill_1 FILLER_99_739 ();
 fill_4 FILLER_99_756 ();
 fill_2 FILLER_99_782 ();
 fill_2 FILLER_99_785 ();
 fill_1 FILLER_99_827 ();
 decap_12 FILLER_99_850 ();
 decap_12 FILLER_99_862 ();
 decap_12 FILLER_99_874 ();
 fill_8 FILLER_99_886 ();
 fill_2 FILLER_99_894 ();
 decap_12 FILLER_99_897 ();
 decap_12 FILLER_99_909 ();
 decap_12 FILLER_99_921 ();
 decap_12 FILLER_99_933 ();
 fill_4 FILLER_99_945 ();
 fill_2 FILLER_99_949 ();
 fill_1 FILLER_99_951 ();
 decap_12 FILLER_99_953 ();
 decap_12 FILLER_99_965 ();
 decap_12 FILLER_99_977 ();
 decap_12 FILLER_99_989 ();
 fill_4 FILLER_99_1001 ();
 fill_2 FILLER_99_1005 ();
 fill_1 FILLER_99_1007 ();
 decap_12 FILLER_99_1009 ();
 decap_12 FILLER_99_1021 ();
 fill_2 FILLER_99_1033 ();
 fill_1 FILLER_100_3 ();
 fill_4 FILLER_100_24 ();
 fill_1 FILLER_100_29 ();
 fill_8 FILLER_100_36 ();
 fill_4 FILLER_100_60 ();
 fill_1 FILLER_100_64 ();
 fill_2 FILLER_100_81 ();
 fill_1 FILLER_100_83 ();
 fill_2 FILLER_100_131 ();
 fill_2 FILLER_100_141 ();
 fill_1 FILLER_100_143 ();
 fill_4 FILLER_100_167 ();
 fill_2 FILLER_100_180 ();
 fill_1 FILLER_100_182 ();
 fill_1 FILLER_100_188 ();
 fill_1 FILLER_100_195 ();
 fill_1 FILLER_100_197 ();
 fill_2 FILLER_100_236 ();
 fill_1 FILLER_100_251 ();
 fill_2 FILLER_100_295 ();
 fill_4 FILLER_100_304 ();
 fill_2 FILLER_100_318 ();
 fill_2 FILLER_100_336 ();
 fill_1 FILLER_100_338 ();
 fill_2 FILLER_100_365 ();
 fill_1 FILLER_100_367 ();
 fill_2 FILLER_100_392 ();
 fill_1 FILLER_100_394 ();
 decap_12 FILLER_100_408 ();
 fill_2 FILLER_100_421 ();
 fill_1 FILLER_100_423 ();
 fill_1 FILLER_100_454 ();
 fill_2 FILLER_100_462 ();
 fill_2 FILLER_100_473 ();
 fill_1 FILLER_100_475 ();
 fill_4 FILLER_100_482 ();
 fill_2 FILLER_100_503 ();
 fill_1 FILLER_100_505 ();
 fill_8 FILLER_100_520 ();
 fill_2 FILLER_100_536 ();
 fill_2 FILLER_100_546 ();
 fill_1 FILLER_100_548 ();
 fill_2 FILLER_100_561 ();
 fill_4 FILLER_100_583 ();
 fill_1 FILLER_100_587 ();
 fill_2 FILLER_100_595 ();
 fill_1 FILLER_100_635 ();
 fill_2 FILLER_100_642 ();
 fill_4 FILLER_100_667 ();
 fill_1 FILLER_100_671 ();
 fill_4 FILLER_100_686 ();
 fill_1 FILLER_100_709 ();
 fill_1 FILLER_100_715 ();
 fill_2 FILLER_100_767 ();
 fill_2 FILLER_100_777 ();
 fill_1 FILLER_100_779 ();
 fill_2 FILLER_100_795 ();
 fill_4 FILLER_100_805 ();
 fill_2 FILLER_100_809 ();
 fill_1 FILLER_100_811 ();
 decap_12 FILLER_100_839 ();
 decap_12 FILLER_100_851 ();
 fill_4 FILLER_100_863 ();
 fill_1 FILLER_100_867 ();
 decap_12 FILLER_100_869 ();
 decap_12 FILLER_100_881 ();
 decap_12 FILLER_100_893 ();
 decap_12 FILLER_100_905 ();
 fill_4 FILLER_100_917 ();
 fill_2 FILLER_100_921 ();
 fill_1 FILLER_100_923 ();
 decap_12 FILLER_100_925 ();
 decap_12 FILLER_100_937 ();
 decap_12 FILLER_100_949 ();
 decap_12 FILLER_100_961 ();
 fill_4 FILLER_100_973 ();
 fill_2 FILLER_100_977 ();
 fill_1 FILLER_100_979 ();
 decap_12 FILLER_100_981 ();
 decap_12 FILLER_100_993 ();
 decap_12 FILLER_100_1005 ();
 decap_12 FILLER_100_1017 ();
 fill_4 FILLER_100_1029 ();
 fill_2 FILLER_100_1033 ();
 fill_1 FILLER_100_1035 ();
 fill_1 FILLER_100_1037 ();
 fill_2 FILLER_101_3 ();
 fill_1 FILLER_101_5 ();
 fill_2 FILLER_101_16 ();
 fill_1 FILLER_101_18 ();
 fill_4 FILLER_101_33 ();
 fill_2 FILLER_101_37 ();
 fill_1 FILLER_101_55 ();
 fill_2 FILLER_101_57 ();
 fill_1 FILLER_101_59 ();
 fill_2 FILLER_101_85 ();
 fill_1 FILLER_101_87 ();
 fill_1 FILLER_101_95 ();
 fill_4 FILLER_101_113 ();
 fill_1 FILLER_101_117 ();
 fill_2 FILLER_101_125 ();
 fill_1 FILLER_101_127 ();
 fill_4 FILLER_101_144 ();
 fill_2 FILLER_101_166 ();
 fill_1 FILLER_101_190 ();
 fill_1 FILLER_101_195 ();
 fill_2 FILLER_101_278 ();
 fill_2 FILLER_101_281 ();
 fill_2 FILLER_101_295 ();
 fill_2 FILLER_101_313 ();
 fill_1 FILLER_101_315 ();
 fill_4 FILLER_101_332 ();
 fill_2 FILLER_101_369 ();
 fill_1 FILLER_101_371 ();
 fill_8 FILLER_101_379 ();
 fill_4 FILLER_101_393 ();
 fill_1 FILLER_101_397 ();
 fill_2 FILLER_101_423 ();
 fill_1 FILLER_101_425 ();
 fill_2 FILLER_101_446 ();
 fill_2 FILLER_101_455 ();
 fill_2 FILLER_101_483 ();
 fill_4 FILLER_101_493 ();
 fill_2 FILLER_101_505 ();
 fill_1 FILLER_101_507 ();
 fill_2 FILLER_101_538 ();
 fill_4 FILLER_101_561 ();
 fill_1 FILLER_101_565 ();
 fill_1 FILLER_101_575 ();
 fill_2 FILLER_101_592 ();
 fill_2 FILLER_101_614 ();
 fill_2 FILLER_101_625 ();
 fill_1 FILLER_101_627 ();
 fill_1 FILLER_101_634 ();
 fill_4 FILLER_101_643 ();
 fill_4 FILLER_101_661 ();
 fill_2 FILLER_101_665 ();
 fill_1 FILLER_101_667 ();
 fill_2 FILLER_101_673 ();
 fill_1 FILLER_101_693 ();
 fill_1 FILLER_101_706 ();
 fill_1 FILLER_101_727 ();
 fill_1 FILLER_101_732 ();
 fill_1 FILLER_101_753 ();
 fill_4 FILLER_101_760 ();
 fill_4 FILLER_101_778 ();
 fill_2 FILLER_101_782 ();
 fill_1 FILLER_101_785 ();
 fill_2 FILLER_101_794 ();
 fill_1 FILLER_101_796 ();
 fill_2 FILLER_101_826 ();
 decap_12 FILLER_101_841 ();
 decap_12 FILLER_101_853 ();
 decap_12 FILLER_101_865 ();
 decap_12 FILLER_101_877 ();
 fill_4 FILLER_101_889 ();
 fill_2 FILLER_101_893 ();
 fill_1 FILLER_101_895 ();
 decap_12 FILLER_101_897 ();
 decap_12 FILLER_101_909 ();
 decap_12 FILLER_101_921 ();
 decap_12 FILLER_101_933 ();
 fill_4 FILLER_101_945 ();
 fill_2 FILLER_101_949 ();
 fill_1 FILLER_101_951 ();
 decap_12 FILLER_101_953 ();
 decap_12 FILLER_101_965 ();
 decap_12 FILLER_101_977 ();
 decap_12 FILLER_101_989 ();
 fill_4 FILLER_101_1001 ();
 fill_2 FILLER_101_1005 ();
 fill_1 FILLER_101_1007 ();
 decap_12 FILLER_101_1009 ();
 decap_12 FILLER_101_1021 ();
 fill_4 FILLER_101_1033 ();
 fill_1 FILLER_101_1037 ();
 fill_1 FILLER_102_3 ();
 fill_1 FILLER_102_27 ();
 fill_4 FILLER_102_29 ();
 fill_2 FILLER_102_33 ();
 fill_1 FILLER_102_35 ();
 fill_2 FILLER_102_85 ();
 fill_1 FILLER_102_103 ();
 fill_4 FILLER_102_127 ();
 fill_2 FILLER_102_138 ();
 fill_2 FILLER_102_147 ();
 fill_1 FILLER_102_149 ();
 fill_1 FILLER_102_171 ();
 fill_1 FILLER_102_179 ();
 fill_2 FILLER_102_188 ();
 fill_2 FILLER_102_246 ();
 fill_1 FILLER_102_278 ();
 fill_1 FILLER_102_292 ();
 fill_4 FILLER_102_316 ();
 fill_1 FILLER_102_345 ();
 fill_2 FILLER_102_362 ();
 fill_1 FILLER_102_385 ();
 fill_1 FILLER_102_396 ();
 fill_2 FILLER_102_411 ();
 fill_2 FILLER_102_421 ();
 fill_1 FILLER_102_430 ();
 fill_4 FILLER_102_457 ();
 fill_2 FILLER_102_461 ();
 fill_1 FILLER_102_471 ();
 fill_2 FILLER_102_487 ();
 fill_1 FILLER_102_489 ();
 fill_1 FILLER_102_522 ();
 fill_1 FILLER_102_531 ();
 fill_1 FILLER_102_553 ();
 fill_4 FILLER_102_560 ();
 fill_1 FILLER_102_564 ();
 fill_2 FILLER_102_585 ();
 fill_1 FILLER_102_587 ();
 fill_1 FILLER_102_593 ();
 fill_8 FILLER_102_601 ();
 fill_2 FILLER_102_609 ();
 fill_1 FILLER_102_614 ();
 fill_2 FILLER_102_623 ();
 fill_8 FILLER_102_636 ();
 fill_4 FILLER_102_653 ();
 fill_1 FILLER_102_657 ();
 fill_2 FILLER_102_668 ();
 fill_4 FILLER_102_682 ();
 fill_1 FILLER_102_699 ();
 fill_1 FILLER_102_709 ();
 fill_1 FILLER_102_726 ();
 fill_2 FILLER_102_747 ();
 fill_4 FILLER_102_793 ();
 fill_1 FILLER_102_797 ();
 decap_12 FILLER_102_847 ();
 fill_8 FILLER_102_859 ();
 fill_1 FILLER_102_867 ();
 decap_12 FILLER_102_869 ();
 decap_12 FILLER_102_881 ();
 decap_12 FILLER_102_893 ();
 decap_12 FILLER_102_905 ();
 fill_4 FILLER_102_917 ();
 fill_2 FILLER_102_921 ();
 fill_1 FILLER_102_923 ();
 decap_12 FILLER_102_925 ();
 decap_12 FILLER_102_937 ();
 decap_12 FILLER_102_949 ();
 decap_12 FILLER_102_961 ();
 fill_4 FILLER_102_973 ();
 fill_2 FILLER_102_977 ();
 fill_1 FILLER_102_979 ();
 decap_12 FILLER_102_981 ();
 decap_12 FILLER_102_993 ();
 decap_12 FILLER_102_1005 ();
 decap_12 FILLER_102_1017 ();
 fill_4 FILLER_102_1029 ();
 fill_2 FILLER_102_1033 ();
 fill_1 FILLER_102_1035 ();
 fill_1 FILLER_102_1037 ();
 decap_12 FILLER_103_3 ();
 fill_2 FILLER_103_15 ();
 fill_1 FILLER_103_17 ();
 fill_4 FILLER_103_89 ();
 fill_1 FILLER_103_93 ();
 fill_4 FILLER_103_113 ();
 fill_2 FILLER_103_117 ();
 fill_1 FILLER_103_119 ();
 fill_1 FILLER_103_129 ();
 fill_4 FILLER_103_146 ();
 fill_2 FILLER_103_150 ();
 fill_1 FILLER_103_169 ();
 fill_2 FILLER_103_221 ();
 fill_1 FILLER_103_223 ();
 fill_1 FILLER_103_225 ();
 fill_1 FILLER_103_242 ();
 fill_2 FILLER_103_250 ();
 fill_1 FILLER_103_272 ();
 fill_2 FILLER_103_281 ();
 fill_2 FILLER_103_346 ();
 fill_1 FILLER_103_391 ();
 fill_1 FILLER_103_420 ();
 fill_4 FILLER_103_441 ();
 fill_1 FILLER_103_449 ();
 fill_2 FILLER_103_453 ();
 fill_2 FILLER_103_465 ();
 fill_4 FILLER_103_474 ();
 fill_4 FILLER_103_488 ();
 fill_2 FILLER_103_508 ();
 fill_1 FILLER_103_510 ();
 fill_1 FILLER_103_516 ();
 fill_1 FILLER_103_520 ();
 fill_1 FILLER_103_540 ();
 fill_2 FILLER_103_547 ();
 fill_1 FILLER_103_549 ();
 fill_2 FILLER_103_581 ();
 fill_2 FILLER_103_604 ();
 fill_2 FILLER_103_614 ();
 fill_2 FILLER_103_632 ();
 fill_2 FILLER_103_648 ();
 fill_1 FILLER_103_650 ();
 fill_1 FILLER_103_667 ();
 fill_1 FILLER_103_696 ();
 fill_2 FILLER_103_717 ();
 fill_2 FILLER_103_726 ();
 fill_2 FILLER_103_781 ();
 fill_1 FILLER_103_783 ();
 fill_1 FILLER_103_795 ();
 fill_2 FILLER_103_802 ();
 fill_8 FILLER_103_824 ();
 fill_1 FILLER_103_839 ();
 decap_12 FILLER_103_841 ();
 decap_12 FILLER_103_853 ();
 decap_12 FILLER_103_865 ();
 decap_12 FILLER_103_877 ();
 fill_4 FILLER_103_889 ();
 fill_2 FILLER_103_893 ();
 fill_1 FILLER_103_895 ();
 decap_12 FILLER_103_897 ();
 decap_12 FILLER_103_909 ();
 decap_12 FILLER_103_921 ();
 decap_12 FILLER_103_933 ();
 fill_4 FILLER_103_945 ();
 fill_2 FILLER_103_949 ();
 fill_1 FILLER_103_951 ();
 decap_12 FILLER_103_953 ();
 decap_12 FILLER_103_965 ();
 decap_12 FILLER_103_977 ();
 decap_12 FILLER_103_989 ();
 fill_4 FILLER_103_1001 ();
 fill_2 FILLER_103_1005 ();
 fill_1 FILLER_103_1007 ();
 decap_12 FILLER_103_1009 ();
 decap_12 FILLER_103_1021 ();
 fill_4 FILLER_103_1033 ();
 fill_1 FILLER_103_1037 ();
 fill_8 FILLER_104_20 ();
 fill_4 FILLER_104_29 ();
 fill_2 FILLER_104_33 ();
 fill_1 FILLER_104_35 ();
 fill_1 FILLER_104_59 ();
 fill_1 FILLER_104_83 ();
 fill_4 FILLER_104_103 ();
 fill_2 FILLER_104_107 ();
 fill_4 FILLER_104_134 ();
 fill_2 FILLER_104_138 ();
 fill_2 FILLER_104_194 ();
 fill_4 FILLER_104_248 ();
 fill_1 FILLER_104_253 ();
 fill_1 FILLER_104_274 ();
 fill_1 FILLER_104_283 ();
 fill_1 FILLER_104_343 ();
 fill_2 FILLER_104_351 ();
 fill_2 FILLER_104_362 ();
 fill_1 FILLER_104_365 ();
 fill_1 FILLER_104_375 ();
 fill_2 FILLER_104_392 ();
 fill_4 FILLER_104_421 ();
 fill_2 FILLER_104_425 ();
 fill_1 FILLER_104_427 ();
 fill_1 FILLER_104_439 ();
 fill_1 FILLER_104_475 ();
 fill_2 FILLER_104_504 ();
 fill_8 FILLER_104_553 ();
 fill_1 FILLER_104_561 ();
 fill_2 FILLER_104_585 ();
 fill_1 FILLER_104_587 ();
 fill_2 FILLER_104_596 ();
 fill_2 FILLER_104_605 ();
 fill_1 FILLER_104_607 ();
 fill_2 FILLER_104_611 ();
 fill_1 FILLER_104_613 ();
 fill_4 FILLER_104_621 ();
 fill_2 FILLER_104_625 ();
 fill_4 FILLER_104_636 ();
 fill_4 FILLER_104_645 ();
 fill_1 FILLER_104_649 ();
 fill_4 FILLER_104_658 ();
 fill_4 FILLER_104_669 ();
 fill_2 FILLER_104_673 ();
 fill_1 FILLER_104_675 ();
 fill_1 FILLER_104_699 ();
 fill_1 FILLER_104_755 ();
 fill_2 FILLER_104_780 ();
 fill_2 FILLER_104_805 ();
 fill_1 FILLER_104_807 ();
 fill_1 FILLER_104_811 ();
 fill_2 FILLER_104_813 ();
 fill_1 FILLER_104_815 ();
 fill_1 FILLER_104_831 ();
 fill_1 FILLER_104_839 ();
 decap_12 FILLER_104_847 ();
 fill_8 FILLER_104_859 ();
 fill_1 FILLER_104_867 ();
 decap_12 FILLER_104_869 ();
 decap_12 FILLER_104_881 ();
 decap_12 FILLER_104_893 ();
 decap_12 FILLER_104_905 ();
 fill_4 FILLER_104_917 ();
 fill_2 FILLER_104_921 ();
 fill_1 FILLER_104_923 ();
 decap_12 FILLER_104_925 ();
 decap_12 FILLER_104_937 ();
 decap_12 FILLER_104_949 ();
 decap_12 FILLER_104_961 ();
 fill_4 FILLER_104_973 ();
 fill_2 FILLER_104_977 ();
 fill_1 FILLER_104_979 ();
 decap_12 FILLER_104_981 ();
 decap_12 FILLER_104_993 ();
 decap_12 FILLER_104_1005 ();
 decap_12 FILLER_104_1017 ();
 fill_4 FILLER_104_1029 ();
 fill_2 FILLER_104_1033 ();
 fill_1 FILLER_104_1035 ();
 fill_1 FILLER_104_1037 ();
 fill_4 FILLER_105_3 ();
 fill_1 FILLER_105_7 ();
 fill_4 FILLER_105_40 ();
 fill_2 FILLER_105_44 ();
 fill_1 FILLER_105_46 ();
 fill_2 FILLER_105_57 ();
 fill_1 FILLER_105_59 ();
 fill_4 FILLER_105_113 ();
 fill_4 FILLER_105_137 ();
 fill_1 FILLER_105_141 ();
 fill_2 FILLER_105_149 ();
 fill_1 FILLER_105_151 ();
 fill_2 FILLER_105_225 ();
 fill_1 FILLER_105_242 ();
 fill_4 FILLER_105_251 ();
 fill_4 FILLER_105_264 ();
 fill_1 FILLER_105_268 ();
 fill_4 FILLER_105_323 ();
 fill_1 FILLER_105_391 ();
 fill_1 FILLER_105_393 ();
 fill_8 FILLER_105_412 ();
 fill_2 FILLER_105_420 ();
 fill_1 FILLER_105_422 ();
 fill_4 FILLER_105_426 ();
 fill_2 FILLER_105_430 ();
 fill_2 FILLER_105_472 ();
 fill_1 FILLER_105_486 ();
 fill_4 FILLER_105_546 ();
 fill_1 FILLER_105_559 ();
 fill_1 FILLER_105_592 ();
 fill_2 FILLER_105_602 ();
 fill_1 FILLER_105_609 ();
 fill_2 FILLER_105_617 ();
 fill_1 FILLER_105_632 ();
 fill_1 FILLER_105_645 ();
 fill_4 FILLER_105_655 ();
 fill_1 FILLER_105_659 ();
 fill_4 FILLER_105_700 ();
 fill_1 FILLER_105_727 ();
 fill_2 FILLER_105_740 ();
 fill_4 FILLER_105_752 ();
 fill_2 FILLER_105_756 ();
 fill_1 FILLER_105_758 ();
 fill_1 FILLER_105_768 ();
 fill_1 FILLER_105_775 ();
 fill_1 FILLER_105_783 ();
 fill_4 FILLER_105_809 ();
 fill_1 FILLER_105_813 ();
 decap_12 FILLER_105_858 ();
 decap_12 FILLER_105_870 ();
 decap_12 FILLER_105_882 ();
 fill_2 FILLER_105_894 ();
 decap_12 FILLER_105_897 ();
 decap_12 FILLER_105_909 ();
 decap_12 FILLER_105_921 ();
 decap_12 FILLER_105_933 ();
 fill_4 FILLER_105_945 ();
 fill_2 FILLER_105_949 ();
 fill_1 FILLER_105_951 ();
 decap_12 FILLER_105_953 ();
 decap_12 FILLER_105_965 ();
 decap_12 FILLER_105_977 ();
 decap_12 FILLER_105_989 ();
 fill_4 FILLER_105_1001 ();
 fill_2 FILLER_105_1005 ();
 fill_1 FILLER_105_1007 ();
 decap_12 FILLER_105_1009 ();
 decap_12 FILLER_105_1021 ();
 fill_4 FILLER_105_1033 ();
 fill_1 FILLER_105_1037 ();
 fill_4 FILLER_106_3 ();
 fill_1 FILLER_106_7 ();
 fill_4 FILLER_106_24 ();
 fill_2 FILLER_106_34 ();
 fill_1 FILLER_106_52 ();
 fill_4 FILLER_106_62 ();
 fill_1 FILLER_106_66 ();
 fill_1 FILLER_106_83 ();
 fill_4 FILLER_106_101 ();
 fill_2 FILLER_106_105 ();
 fill_1 FILLER_106_107 ();
 fill_2 FILLER_106_115 ();
 fill_2 FILLER_106_168 ();
 fill_1 FILLER_106_186 ();
 fill_2 FILLER_106_194 ();
 fill_2 FILLER_106_206 ();
 fill_1 FILLER_106_208 ();
 fill_1 FILLER_106_219 ();
 fill_4 FILLER_106_233 ();
 fill_2 FILLER_106_237 ();
 fill_1 FILLER_106_239 ();
 fill_1 FILLER_106_251 ();
 fill_2 FILLER_106_253 ();
 fill_2 FILLER_106_262 ();
 fill_1 FILLER_106_273 ();
 fill_2 FILLER_106_277 ();
 fill_1 FILLER_106_365 ();
 fill_1 FILLER_106_395 ();
 fill_2 FILLER_106_417 ();
 fill_1 FILLER_106_419 ();
 fill_2 FILLER_106_452 ();
 fill_2 FILLER_106_474 ();
 fill_1 FILLER_106_485 ();
 fill_1 FILLER_106_503 ();
 fill_2 FILLER_106_517 ();
 fill_1 FILLER_106_531 ();
 fill_8 FILLER_106_533 ();
 fill_1 FILLER_106_541 ();
 fill_2 FILLER_106_550 ();
 fill_1 FILLER_106_552 ();
 fill_4 FILLER_106_565 ();
 fill_8 FILLER_106_578 ();
 fill_2 FILLER_106_586 ();
 fill_2 FILLER_106_617 ();
 fill_2 FILLER_106_642 ();
 fill_8 FILLER_106_668 ();
 fill_1 FILLER_106_676 ();
 fill_4 FILLER_106_680 ();
 fill_4 FILLER_106_691 ();
 fill_2 FILLER_106_695 ();
 fill_2 FILLER_106_760 ();
 fill_1 FILLER_106_762 ();
 fill_4 FILLER_106_790 ();
 fill_8 FILLER_106_802 ();
 fill_2 FILLER_106_810 ();
 fill_4 FILLER_106_827 ();
 fill_2 FILLER_106_835 ();
 decap_12 FILLER_106_840 ();
 decap_12 FILLER_106_852 ();
 fill_4 FILLER_106_864 ();
 decap_12 FILLER_106_869 ();
 decap_12 FILLER_106_881 ();
 decap_12 FILLER_106_893 ();
 decap_12 FILLER_106_905 ();
 fill_4 FILLER_106_917 ();
 fill_2 FILLER_106_921 ();
 fill_1 FILLER_106_923 ();
 decap_12 FILLER_106_925 ();
 decap_12 FILLER_106_937 ();
 decap_12 FILLER_106_949 ();
 decap_12 FILLER_106_961 ();
 fill_4 FILLER_106_973 ();
 fill_2 FILLER_106_977 ();
 fill_1 FILLER_106_979 ();
 decap_12 FILLER_106_981 ();
 decap_12 FILLER_106_993 ();
 decap_12 FILLER_106_1005 ();
 decap_12 FILLER_106_1017 ();
 fill_4 FILLER_106_1029 ();
 fill_2 FILLER_106_1033 ();
 fill_1 FILLER_106_1035 ();
 fill_1 FILLER_106_1037 ();
 fill_2 FILLER_107_38 ();
 fill_1 FILLER_107_64 ();
 fill_4 FILLER_107_169 ();
 fill_2 FILLER_107_218 ();
 fill_4 FILLER_107_300 ();
 fill_2 FILLER_107_304 ();
 fill_1 FILLER_107_306 ();
 fill_2 FILLER_107_351 ();
 fill_1 FILLER_107_353 ();
 fill_1 FILLER_107_399 ();
 fill_2 FILLER_107_423 ();
 fill_2 FILLER_107_432 ();
 fill_2 FILLER_107_455 ();
 fill_1 FILLER_107_477 ();
 fill_1 FILLER_107_503 ();
 fill_2 FILLER_107_541 ();
 fill_1 FILLER_107_543 ();
 fill_2 FILLER_107_553 ();
 fill_1 FILLER_107_555 ();
 fill_1 FILLER_107_559 ();
 fill_2 FILLER_107_588 ();
 fill_4 FILLER_107_593 ();
 fill_1 FILLER_107_603 ();
 fill_1 FILLER_107_615 ();
 fill_1 FILLER_107_621 ();
 fill_4 FILLER_107_638 ();
 fill_2 FILLER_107_642 ();
 fill_2 FILLER_107_647 ();
 fill_1 FILLER_107_649 ();
 fill_2 FILLER_107_673 ();
 fill_4 FILLER_107_695 ();
 fill_1 FILLER_107_699 ();
 fill_2 FILLER_107_703 ();
 fill_2 FILLER_107_737 ();
 fill_2 FILLER_107_752 ();
 fill_4 FILLER_107_766 ();
 fill_4 FILLER_107_779 ();
 fill_1 FILLER_107_783 ();
 fill_2 FILLER_107_785 ();
 fill_1 FILLER_107_787 ();
 fill_2 FILLER_107_816 ();
 fill_1 FILLER_107_818 ();
 fill_2 FILLER_107_826 ();
 fill_1 FILLER_107_828 ();
 fill_4 FILLER_107_834 ();
 fill_2 FILLER_107_838 ();
 decap_12 FILLER_107_848 ();
 decap_12 FILLER_107_860 ();
 decap_12 FILLER_107_872 ();
 decap_12 FILLER_107_884 ();
 decap_12 FILLER_107_897 ();
 decap_12 FILLER_107_909 ();
 decap_12 FILLER_107_921 ();
 decap_12 FILLER_107_933 ();
 fill_4 FILLER_107_945 ();
 fill_2 FILLER_107_949 ();
 fill_1 FILLER_107_951 ();
 decap_12 FILLER_107_953 ();
 decap_12 FILLER_107_965 ();
 decap_12 FILLER_107_977 ();
 decap_12 FILLER_107_989 ();
 fill_4 FILLER_107_1001 ();
 fill_2 FILLER_107_1005 ();
 fill_1 FILLER_107_1007 ();
 decap_12 FILLER_107_1009 ();
 decap_12 FILLER_107_1021 ();
 fill_4 FILLER_107_1033 ();
 fill_1 FILLER_107_1037 ();
 fill_2 FILLER_108_3 ();
 fill_4 FILLER_108_21 ();
 fill_2 FILLER_108_25 ();
 fill_1 FILLER_108_27 ();
 fill_2 FILLER_108_35 ();
 fill_1 FILLER_108_37 ();
 fill_8 FILLER_108_45 ();
 fill_2 FILLER_108_53 ();
 fill_1 FILLER_108_55 ();
 fill_1 FILLER_108_99 ();
 fill_2 FILLER_108_123 ();
 fill_1 FILLER_108_125 ();
 fill_1 FILLER_108_145 ();
 fill_1 FILLER_108_158 ();
 fill_2 FILLER_108_194 ();
 fill_2 FILLER_108_210 ();
 fill_2 FILLER_108_219 ();
 fill_1 FILLER_108_221 ();
 fill_8 FILLER_108_229 ();
 fill_1 FILLER_108_237 ();
 fill_2 FILLER_108_253 ();
 fill_1 FILLER_108_255 ();
 fill_4 FILLER_108_276 ();
 fill_2 FILLER_108_280 ();
 fill_2 FILLER_108_306 ();
 fill_4 FILLER_108_309 ();
 fill_2 FILLER_108_313 ();
 fill_1 FILLER_108_359 ();
 fill_1 FILLER_108_421 ();
 fill_2 FILLER_108_442 ();
 fill_1 FILLER_108_463 ();
 fill_1 FILLER_108_533 ();
 fill_4 FILLER_108_542 ();
 fill_1 FILLER_108_555 ();
 fill_8 FILLER_108_562 ();
 fill_1 FILLER_108_580 ();
 fill_1 FILLER_108_587 ();
 fill_1 FILLER_108_603 ();
 fill_2 FILLER_108_614 ();
 fill_1 FILLER_108_623 ();
 fill_1 FILLER_108_662 ();
 fill_1 FILLER_108_692 ();
 fill_2 FILLER_108_698 ();
 decap_12 FILLER_108_701 ();
 fill_2 FILLER_108_713 ();
 fill_1 FILLER_108_715 ();
 fill_4 FILLER_108_723 ();
 fill_2 FILLER_108_727 ();
 fill_1 FILLER_108_729 ();
 fill_1 FILLER_108_757 ();
 fill_1 FILLER_108_765 ();
 fill_1 FILLER_108_779 ();
 fill_4 FILLER_108_793 ();
 fill_2 FILLER_108_800 ();
 fill_1 FILLER_108_802 ();
 fill_2 FILLER_108_818 ();
 fill_2 FILLER_108_826 ();
 fill_1 FILLER_108_828 ();
 decap_12 FILLER_108_847 ();
 fill_8 FILLER_108_859 ();
 fill_1 FILLER_108_867 ();
 decap_12 FILLER_108_869 ();
 decap_12 FILLER_108_881 ();
 decap_12 FILLER_108_893 ();
 decap_12 FILLER_108_905 ();
 fill_4 FILLER_108_917 ();
 fill_2 FILLER_108_921 ();
 fill_1 FILLER_108_923 ();
 decap_12 FILLER_108_925 ();
 decap_12 FILLER_108_937 ();
 decap_12 FILLER_108_949 ();
 decap_12 FILLER_108_961 ();
 fill_4 FILLER_108_973 ();
 fill_2 FILLER_108_977 ();
 fill_1 FILLER_108_979 ();
 decap_12 FILLER_108_981 ();
 decap_12 FILLER_108_993 ();
 decap_12 FILLER_108_1005 ();
 fill_8 FILLER_108_1017 ();
 fill_1 FILLER_108_1025 ();
 fill_1 FILLER_108_1037 ();
 fill_1 FILLER_109_19 ();
 fill_1 FILLER_109_55 ();
 fill_2 FILLER_109_86 ();
 fill_1 FILLER_109_88 ();
 fill_4 FILLER_109_97 ();
 fill_1 FILLER_109_101 ();
 fill_2 FILLER_109_110 ();
 fill_1 FILLER_109_121 ();
 fill_2 FILLER_109_146 ();
 fill_1 FILLER_109_161 ();
 fill_2 FILLER_109_165 ();
 fill_1 FILLER_109_167 ();
 fill_4 FILLER_109_178 ();
 fill_2 FILLER_109_182 ();
 fill_2 FILLER_109_245 ();
 fill_2 FILLER_109_284 ();
 fill_1 FILLER_109_290 ();
 fill_2 FILLER_109_320 ();
 fill_1 FILLER_109_322 ();
 fill_2 FILLER_109_337 ();
 fill_4 FILLER_109_409 ();
 fill_1 FILLER_109_413 ();
 fill_2 FILLER_109_420 ();
 fill_1 FILLER_109_422 ();
 fill_1 FILLER_109_426 ();
 fill_1 FILLER_109_477 ();
 fill_2 FILLER_109_510 ();
 fill_4 FILLER_109_549 ();
 fill_1 FILLER_109_591 ();
 fill_1 FILLER_109_595 ();
 fill_1 FILLER_109_604 ();
 fill_2 FILLER_109_653 ();
 fill_1 FILLER_109_655 ();
 fill_4 FILLER_109_667 ();
 fill_1 FILLER_109_671 ();
 fill_8 FILLER_109_673 ();
 fill_2 FILLER_109_681 ();
 fill_2 FILLER_109_688 ();
 fill_1 FILLER_109_690 ();
 fill_1 FILLER_109_720 ();
 fill_2 FILLER_109_766 ();
 fill_2 FILLER_109_774 ();
 fill_1 FILLER_109_790 ();
 fill_2 FILLER_109_806 ();
 fill_1 FILLER_109_808 ();
 fill_2 FILLER_109_812 ();
 fill_1 FILLER_109_818 ();
 fill_4 FILLER_109_824 ();
 fill_2 FILLER_109_828 ();
 fill_1 FILLER_109_830 ();
 decap_12 FILLER_109_846 ();
 decap_12 FILLER_109_858 ();
 decap_12 FILLER_109_870 ();
 decap_12 FILLER_109_882 ();
 fill_2 FILLER_109_894 ();
 decap_12 FILLER_109_897 ();
 decap_12 FILLER_109_909 ();
 decap_12 FILLER_109_921 ();
 decap_12 FILLER_109_933 ();
 fill_4 FILLER_109_945 ();
 fill_2 FILLER_109_949 ();
 fill_1 FILLER_109_951 ();
 decap_12 FILLER_109_953 ();
 decap_12 FILLER_109_965 ();
 decap_12 FILLER_109_977 ();
 decap_12 FILLER_109_989 ();
 fill_4 FILLER_109_1001 ();
 fill_2 FILLER_109_1005 ();
 fill_1 FILLER_109_1007 ();
 decap_12 FILLER_109_1009 ();
 decap_12 FILLER_109_1021 ();
 fill_4 FILLER_109_1033 ();
 fill_1 FILLER_109_1037 ();
 decap_12 FILLER_110_3 ();
 fill_2 FILLER_110_20 ();
 fill_1 FILLER_110_22 ();
 fill_2 FILLER_110_26 ();
 fill_1 FILLER_110_32 ();
 fill_1 FILLER_110_38 ();
 fill_2 FILLER_110_48 ();
 fill_4 FILLER_110_85 ();
 fill_2 FILLER_110_89 ();
 fill_1 FILLER_110_91 ();
 fill_1 FILLER_110_116 ();
 fill_4 FILLER_110_134 ();
 fill_2 FILLER_110_138 ();
 fill_2 FILLER_110_141 ();
 fill_1 FILLER_110_143 ();
 fill_2 FILLER_110_152 ();
 fill_4 FILLER_110_168 ();
 fill_1 FILLER_110_206 ();
 fill_4 FILLER_110_225 ();
 fill_1 FILLER_110_229 ();
 fill_2 FILLER_110_250 ();
 fill_2 FILLER_110_265 ();
 fill_2 FILLER_110_276 ();
 fill_1 FILLER_110_301 ();
 fill_1 FILLER_110_357 ();
 fill_1 FILLER_110_373 ();
 fill_1 FILLER_110_437 ();
 fill_2 FILLER_110_450 ();
 fill_1 FILLER_110_531 ();
 fill_1 FILLER_110_537 ();
 fill_4 FILLER_110_554 ();
 fill_2 FILLER_110_558 ();
 fill_8 FILLER_110_565 ();
 fill_2 FILLER_110_576 ();
 fill_1 FILLER_110_578 ();
 fill_4 FILLER_110_582 ();
 fill_2 FILLER_110_586 ();
 fill_4 FILLER_110_589 ();
 fill_8 FILLER_110_599 ();
 fill_2 FILLER_110_607 ();
 fill_4 FILLER_110_625 ();
 fill_4 FILLER_110_638 ();
 fill_2 FILLER_110_642 ();
 fill_2 FILLER_110_668 ();
 fill_1 FILLER_110_670 ();
 fill_8 FILLER_110_692 ();
 fill_2 FILLER_110_701 ();
 fill_1 FILLER_110_703 ();
 fill_4 FILLER_110_727 ();
 fill_2 FILLER_110_738 ();
 fill_4 FILLER_110_757 ();
 fill_2 FILLER_110_796 ();
 fill_1 FILLER_110_798 ();
 fill_4 FILLER_110_802 ();
 fill_1 FILLER_110_829 ();
 fill_1 FILLER_110_844 ();
 fill_2 FILLER_110_865 ();
 fill_1 FILLER_110_867 ();
 decap_12 FILLER_110_877 ();
 decap_12 FILLER_110_889 ();
 decap_12 FILLER_110_901 ();
 fill_8 FILLER_110_913 ();
 fill_2 FILLER_110_921 ();
 fill_1 FILLER_110_923 ();
 decap_12 FILLER_110_925 ();
 decap_12 FILLER_110_937 ();
 decap_12 FILLER_110_949 ();
 decap_12 FILLER_110_961 ();
 fill_4 FILLER_110_973 ();
 fill_2 FILLER_110_977 ();
 fill_1 FILLER_110_979 ();
 decap_12 FILLER_110_981 ();
 decap_12 FILLER_110_993 ();
 decap_12 FILLER_110_1005 ();
 decap_12 FILLER_110_1017 ();
 fill_4 FILLER_110_1029 ();
 fill_2 FILLER_110_1033 ();
 fill_1 FILLER_110_1035 ();
 fill_1 FILLER_110_1037 ();
 decap_12 FILLER_111_7 ();
 fill_4 FILLER_111_19 ();
 fill_1 FILLER_111_23 ();
 fill_2 FILLER_111_37 ();
 fill_4 FILLER_111_52 ();
 fill_4 FILLER_111_107 ();
 fill_1 FILLER_111_111 ();
 fill_2 FILLER_111_113 ();
 fill_1 FILLER_111_115 ();
 fill_1 FILLER_111_124 ();
 fill_2 FILLER_111_132 ();
 fill_2 FILLER_111_149 ();
 fill_1 FILLER_111_160 ();
 fill_2 FILLER_111_169 ();
 fill_1 FILLER_111_186 ();
 fill_1 FILLER_111_192 ();
 fill_1 FILLER_111_198 ();
 fill_2 FILLER_111_222 ();
 fill_2 FILLER_111_242 ();
 fill_2 FILLER_111_278 ();
 fill_1 FILLER_111_285 ();
 fill_1 FILLER_111_306 ();
 fill_1 FILLER_111_322 ();
 fill_2 FILLER_111_350 ();
 fill_1 FILLER_111_359 ();
 fill_1 FILLER_111_376 ();
 fill_2 FILLER_111_396 ();
 fill_1 FILLER_111_434 ();
 fill_1 FILLER_111_447 ();
 fill_1 FILLER_111_503 ();
 fill_2 FILLER_111_514 ();
 fill_8 FILLER_111_532 ();
 fill_8 FILLER_111_546 ();
 fill_4 FILLER_111_570 ();
 fill_2 FILLER_111_584 ();
 fill_1 FILLER_111_589 ();
 fill_4 FILLER_111_597 ();
 fill_4 FILLER_111_610 ();
 fill_2 FILLER_111_614 ();
 fill_2 FILLER_111_617 ();
 fill_8 FILLER_111_639 ();
 fill_1 FILLER_111_686 ();
 fill_2 FILLER_111_725 ();
 fill_1 FILLER_111_727 ();
 fill_4 FILLER_111_761 ();
 fill_1 FILLER_111_765 ();
 fill_4 FILLER_111_775 ();
 fill_2 FILLER_111_779 ();
 fill_8 FILLER_111_801 ();
 fill_1 FILLER_111_809 ();
 fill_2 FILLER_111_819 ();
 fill_1 FILLER_111_821 ();
 fill_4 FILLER_111_833 ();
 fill_2 FILLER_111_837 ();
 fill_1 FILLER_111_839 ();
 fill_4 FILLER_111_844 ();
 fill_1 FILLER_111_851 ();
 fill_2 FILLER_111_857 ();
 fill_4 FILLER_111_889 ();
 fill_2 FILLER_111_893 ();
 fill_1 FILLER_111_895 ();
 decap_12 FILLER_111_897 ();
 decap_12 FILLER_111_909 ();
 decap_12 FILLER_111_921 ();
 decap_12 FILLER_111_933 ();
 fill_4 FILLER_111_945 ();
 fill_2 FILLER_111_949 ();
 fill_1 FILLER_111_951 ();
 decap_12 FILLER_111_953 ();
 decap_12 FILLER_111_965 ();
 decap_12 FILLER_111_977 ();
 decap_12 FILLER_111_989 ();
 fill_4 FILLER_111_1001 ();
 fill_2 FILLER_111_1005 ();
 fill_1 FILLER_111_1007 ();
 decap_12 FILLER_111_1009 ();
 decap_12 FILLER_111_1021 ();
 fill_4 FILLER_111_1033 ();
 fill_1 FILLER_111_1037 ();
 decap_12 FILLER_112_3 ();
 decap_12 FILLER_112_15 ();
 fill_1 FILLER_112_27 ();
 fill_1 FILLER_112_45 ();
 fill_2 FILLER_112_71 ();
 fill_2 FILLER_112_81 ();
 fill_1 FILLER_112_83 ();
 fill_2 FILLER_112_85 ();
 fill_1 FILLER_112_90 ();
 fill_4 FILLER_112_99 ();
 fill_1 FILLER_112_103 ();
 fill_1 FILLER_112_130 ();
 fill_2 FILLER_112_151 ();
 fill_2 FILLER_112_158 ();
 fill_1 FILLER_112_176 ();
 fill_2 FILLER_112_188 ();
 fill_1 FILLER_112_190 ();
 fill_2 FILLER_112_194 ();
 fill_1 FILLER_112_197 ();
 fill_2 FILLER_112_216 ();
 fill_2 FILLER_112_253 ();
 fill_1 FILLER_112_255 ();
 fill_2 FILLER_112_263 ();
 fill_1 FILLER_112_265 ();
 fill_2 FILLER_112_286 ();
 fill_2 FILLER_112_298 ();
 fill_1 FILLER_112_309 ();
 fill_1 FILLER_112_324 ();
 fill_2 FILLER_112_332 ();
 fill_1 FILLER_112_357 ();
 fill_2 FILLER_112_365 ();
 fill_1 FILLER_112_389 ();
 fill_2 FILLER_112_410 ();
 fill_2 FILLER_112_464 ();
 fill_2 FILLER_112_477 ();
 fill_1 FILLER_112_531 ();
 fill_2 FILLER_112_546 ();
 fill_1 FILLER_112_548 ();
 fill_2 FILLER_112_557 ();
 fill_1 FILLER_112_559 ();
 fill_2 FILLER_112_586 ();
 decap_12 FILLER_112_630 ();
 fill_2 FILLER_112_642 ();
 fill_2 FILLER_112_659 ();
 fill_8 FILLER_112_689 ();
 fill_2 FILLER_112_697 ();
 fill_1 FILLER_112_699 ();
 fill_1 FILLER_112_737 ();
 fill_2 FILLER_112_741 ();
 fill_2 FILLER_112_746 ();
 fill_1 FILLER_112_748 ();
 fill_4 FILLER_112_752 ();
 fill_8 FILLER_112_781 ();
 fill_2 FILLER_112_801 ();
 fill_8 FILLER_112_829 ();
 fill_4 FILLER_112_863 ();
 fill_1 FILLER_112_867 ();
 decap_12 FILLER_112_889 ();
 decap_12 FILLER_112_901 ();
 fill_8 FILLER_112_913 ();
 fill_2 FILLER_112_921 ();
 fill_1 FILLER_112_923 ();
 decap_12 FILLER_112_925 ();
 decap_12 FILLER_112_937 ();
 decap_12 FILLER_112_949 ();
 decap_12 FILLER_112_961 ();
 fill_4 FILLER_112_973 ();
 fill_2 FILLER_112_977 ();
 fill_1 FILLER_112_979 ();
 decap_12 FILLER_112_981 ();
 decap_12 FILLER_112_993 ();
 decap_12 FILLER_112_1005 ();
 decap_12 FILLER_112_1017 ();
 fill_4 FILLER_112_1029 ();
 fill_2 FILLER_112_1033 ();
 fill_1 FILLER_112_1035 ();
 fill_1 FILLER_112_1037 ();
 decap_12 FILLER_113_3 ();
 decap_12 FILLER_113_15 ();
 fill_1 FILLER_113_55 ();
 fill_4 FILLER_113_61 ();
 fill_1 FILLER_113_65 ();
 fill_2 FILLER_113_109 ();
 fill_1 FILLER_113_111 ();
 fill_1 FILLER_113_177 ();
 fill_2 FILLER_113_208 ();
 fill_1 FILLER_113_225 ();
 fill_4 FILLER_113_271 ();
 fill_2 FILLER_113_275 ();
 fill_1 FILLER_113_335 ();
 fill_1 FILLER_113_348 ();
 fill_1 FILLER_113_366 ();
 fill_2 FILLER_113_390 ();
 fill_2 FILLER_113_406 ();
 fill_1 FILLER_113_436 ();
 fill_4 FILLER_113_452 ();
 fill_1 FILLER_113_456 ();
 fill_2 FILLER_113_470 ();
 fill_2 FILLER_113_489 ();
 fill_1 FILLER_113_513 ();
 fill_4 FILLER_113_547 ();
 fill_2 FILLER_113_551 ();
 fill_1 FILLER_113_553 ();
 fill_2 FILLER_113_557 ();
 fill_1 FILLER_113_559 ();
 decap_12 FILLER_113_573 ();
 fill_1 FILLER_113_598 ();
 fill_1 FILLER_113_641 ();
 fill_1 FILLER_113_652 ();
 fill_4 FILLER_113_667 ();
 fill_1 FILLER_113_671 ();
 fill_2 FILLER_113_673 ();
 fill_2 FILLER_113_679 ();
 fill_2 FILLER_113_690 ();
 fill_4 FILLER_113_721 ();
 fill_2 FILLER_113_725 ();
 fill_1 FILLER_113_727 ();
 fill_2 FILLER_113_750 ();
 fill_1 FILLER_113_771 ();
 fill_1 FILLER_113_783 ();
 fill_1 FILLER_113_839 ();
 fill_2 FILLER_113_893 ();
 fill_1 FILLER_113_895 ();
 decap_12 FILLER_113_897 ();
 decap_12 FILLER_113_909 ();
 decap_12 FILLER_113_921 ();
 decap_12 FILLER_113_933 ();
 fill_4 FILLER_113_945 ();
 fill_2 FILLER_113_949 ();
 fill_1 FILLER_113_951 ();
 decap_12 FILLER_113_953 ();
 decap_12 FILLER_113_965 ();
 decap_12 FILLER_113_977 ();
 decap_12 FILLER_113_989 ();
 fill_4 FILLER_113_1001 ();
 fill_2 FILLER_113_1005 ();
 fill_1 FILLER_113_1007 ();
 decap_12 FILLER_113_1009 ();
 decap_12 FILLER_113_1021 ();
 fill_4 FILLER_113_1033 ();
 fill_1 FILLER_113_1037 ();
 decap_12 FILLER_114_3 ();
 decap_12 FILLER_114_15 ();
 fill_1 FILLER_114_27 ();
 decap_12 FILLER_114_29 ();
 fill_8 FILLER_114_61 ();
 fill_4 FILLER_114_78 ();
 fill_2 FILLER_114_82 ();
 fill_1 FILLER_114_94 ();
 fill_2 FILLER_114_115 ();
 fill_2 FILLER_114_137 ();
 fill_1 FILLER_114_139 ();
 fill_2 FILLER_114_141 ();
 fill_2 FILLER_114_150 ();
 fill_4 FILLER_114_192 ();
 fill_4 FILLER_114_200 ();
 fill_1 FILLER_114_213 ();
 fill_1 FILLER_114_245 ();
 fill_2 FILLER_114_260 ();
 fill_1 FILLER_114_350 ();
 fill_1 FILLER_114_365 ();
 fill_1 FILLER_114_377 ();
 fill_2 FILLER_114_401 ();
 decap_12 FILLER_114_445 ();
 fill_4 FILLER_114_457 ();
 fill_2 FILLER_114_461 ();
 fill_1 FILLER_114_463 ();
 fill_1 FILLER_114_477 ();
 fill_1 FILLER_114_481 ();
 fill_2 FILLER_114_498 ();
 fill_2 FILLER_114_533 ();
 fill_4 FILLER_114_542 ();
 fill_2 FILLER_114_579 ();
 fill_1 FILLER_114_587 ();
 fill_4 FILLER_114_592 ();
 fill_2 FILLER_114_621 ();
 fill_1 FILLER_114_623 ();
 fill_2 FILLER_114_660 ();
 fill_4 FILLER_114_695 ();
 fill_1 FILLER_114_699 ();
 fill_4 FILLER_114_701 ();
 fill_1 FILLER_114_717 ();
 fill_2 FILLER_114_729 ();
 fill_4 FILLER_114_748 ();
 fill_1 FILLER_114_752 ();
 fill_1 FILLER_114_772 ();
 fill_2 FILLER_114_782 ();
 fill_1 FILLER_114_784 ();
 fill_4 FILLER_114_793 ();
 fill_2 FILLER_114_797 ();
 fill_4 FILLER_114_808 ();
 fill_4 FILLER_114_813 ();
 fill_2 FILLER_114_817 ();
 fill_1 FILLER_114_819 ();
 fill_2 FILLER_114_836 ();
 fill_2 FILLER_114_858 ();
 decap_12 FILLER_114_895 ();
 decap_12 FILLER_114_907 ();
 fill_4 FILLER_114_919 ();
 fill_1 FILLER_114_923 ();
 decap_12 FILLER_114_925 ();
 decap_12 FILLER_114_937 ();
 decap_12 FILLER_114_949 ();
 decap_12 FILLER_114_961 ();
 fill_4 FILLER_114_973 ();
 fill_2 FILLER_114_977 ();
 fill_1 FILLER_114_979 ();
 decap_12 FILLER_114_981 ();
 decap_12 FILLER_114_993 ();
 decap_12 FILLER_114_1005 ();
 decap_12 FILLER_114_1017 ();
 fill_4 FILLER_114_1029 ();
 fill_2 FILLER_114_1033 ();
 fill_1 FILLER_114_1035 ();
 fill_1 FILLER_114_1037 ();
 decap_12 FILLER_115_3 ();
 decap_12 FILLER_115_15 ();
 decap_12 FILLER_115_27 ();
 decap_12 FILLER_115_39 ();
 fill_4 FILLER_115_51 ();
 fill_1 FILLER_115_55 ();
 fill_1 FILLER_115_95 ();
 fill_2 FILLER_115_146 ();
 fill_1 FILLER_115_148 ();
 fill_1 FILLER_115_175 ();
 fill_2 FILLER_115_215 ();
 fill_1 FILLER_115_247 ();
 fill_2 FILLER_115_262 ();
 fill_2 FILLER_115_277 ();
 fill_1 FILLER_115_279 ();
 fill_1 FILLER_115_281 ();
 fill_1 FILLER_115_287 ();
 fill_2 FILLER_115_292 ();
 fill_2 FILLER_115_309 ();
 fill_1 FILLER_115_311 ();
 fill_2 FILLER_115_357 ();
 fill_1 FILLER_115_400 ();
 fill_2 FILLER_115_458 ();
 fill_1 FILLER_115_503 ();
 fill_1 FILLER_115_559 ();
 fill_2 FILLER_115_561 ();
 fill_1 FILLER_115_563 ();
 fill_1 FILLER_115_584 ();
 fill_2 FILLER_115_614 ();
 fill_1 FILLER_115_633 ();
 fill_4 FILLER_115_655 ();
 fill_2 FILLER_115_670 ();
 fill_1 FILLER_115_733 ();
 fill_4 FILLER_115_777 ();
 fill_2 FILLER_115_781 ();
 fill_1 FILLER_115_783 ();
 fill_2 FILLER_115_785 ();
 fill_1 FILLER_115_787 ();
 fill_4 FILLER_115_791 ();
 fill_2 FILLER_115_795 ();
 fill_2 FILLER_115_838 ();
 fill_1 FILLER_115_867 ();
 fill_8 FILLER_115_885 ();
 fill_2 FILLER_115_893 ();
 fill_1 FILLER_115_895 ();
 decap_12 FILLER_115_897 ();
 decap_12 FILLER_115_909 ();
 decap_12 FILLER_115_921 ();
 decap_12 FILLER_115_933 ();
 fill_4 FILLER_115_945 ();
 fill_2 FILLER_115_949 ();
 fill_1 FILLER_115_951 ();
 decap_12 FILLER_115_953 ();
 decap_12 FILLER_115_965 ();
 decap_12 FILLER_115_977 ();
 decap_12 FILLER_115_989 ();
 fill_4 FILLER_115_1001 ();
 fill_2 FILLER_115_1005 ();
 fill_1 FILLER_115_1007 ();
 decap_12 FILLER_115_1009 ();
 decap_12 FILLER_115_1021 ();
 fill_4 FILLER_115_1033 ();
 fill_1 FILLER_115_1037 ();
 decap_12 FILLER_116_3 ();
 decap_12 FILLER_116_15 ();
 fill_1 FILLER_116_27 ();
 decap_12 FILLER_116_29 ();
 decap_12 FILLER_116_41 ();
 decap_12 FILLER_116_53 ();
 fill_2 FILLER_116_65 ();
 fill_1 FILLER_116_67 ();
 fill_4 FILLER_116_78 ();
 fill_2 FILLER_116_82 ();
 fill_2 FILLER_116_187 ();
 fill_2 FILLER_116_205 ();
 fill_2 FILLER_116_215 ();
 fill_1 FILLER_116_225 ();
 fill_1 FILLER_116_231 ();
 fill_2 FILLER_116_250 ();
 fill_1 FILLER_116_267 ();
 fill_1 FILLER_116_275 ();
 fill_2 FILLER_116_306 ();
 fill_2 FILLER_116_317 ();
 fill_2 FILLER_116_332 ();
 fill_1 FILLER_116_348 ();
 fill_1 FILLER_116_356 ();
 fill_1 FILLER_116_363 ();
 fill_1 FILLER_116_371 ();
 fill_1 FILLER_116_381 ();
 fill_2 FILLER_116_386 ();
 fill_1 FILLER_116_399 ();
 fill_2 FILLER_116_414 ();
 fill_1 FILLER_116_416 ();
 fill_1 FILLER_116_447 ();
 fill_1 FILLER_116_455 ();
 fill_1 FILLER_116_466 ();
 fill_1 FILLER_116_507 ();
 fill_4 FILLER_116_516 ();
 fill_2 FILLER_116_520 ();
 fill_1 FILLER_116_522 ();
 fill_1 FILLER_116_531 ();
 fill_1 FILLER_116_536 ();
 fill_1 FILLER_116_544 ();
 fill_2 FILLER_116_552 ();
 fill_2 FILLER_116_570 ();
 fill_1 FILLER_116_572 ();
 fill_1 FILLER_116_587 ();
 fill_2 FILLER_116_593 ();
 fill_1 FILLER_116_611 ();
 fill_1 FILLER_116_643 ();
 fill_4 FILLER_116_661 ();
 fill_2 FILLER_116_697 ();
 fill_1 FILLER_116_699 ();
 fill_2 FILLER_116_701 ();
 fill_1 FILLER_116_703 ();
 fill_1 FILLER_116_741 ();
 fill_1 FILLER_116_771 ();
 fill_4 FILLER_116_805 ();
 fill_2 FILLER_116_809 ();
 fill_1 FILLER_116_811 ();
 fill_4 FILLER_116_822 ();
 fill_2 FILLER_116_826 ();
 fill_1 FILLER_116_839 ();
 fill_2 FILLER_116_869 ();
 fill_1 FILLER_116_871 ();
 decap_12 FILLER_116_893 ();
 fill_8 FILLER_116_905 ();
 fill_1 FILLER_116_913 ();
 fill_4 FILLER_116_918 ();
 fill_2 FILLER_116_922 ();
 fill_1 FILLER_116_925 ();
 decap_12 FILLER_116_934 ();
 decap_12 FILLER_116_946 ();
 decap_12 FILLER_116_958 ();
 fill_8 FILLER_116_970 ();
 fill_2 FILLER_116_978 ();
 decap_12 FILLER_116_981 ();
 decap_12 FILLER_116_993 ();
 decap_12 FILLER_116_1005 ();
 decap_12 FILLER_116_1017 ();
 fill_4 FILLER_116_1029 ();
 fill_2 FILLER_116_1033 ();
 fill_1 FILLER_116_1035 ();
 fill_1 FILLER_116_1037 ();
 decap_12 FILLER_117_3 ();
 decap_12 FILLER_117_15 ();
 decap_12 FILLER_117_27 ();
 decap_12 FILLER_117_39 ();
 fill_4 FILLER_117_51 ();
 fill_1 FILLER_117_55 ();
 fill_8 FILLER_117_57 ();
 fill_2 FILLER_117_65 ();
 fill_8 FILLER_117_76 ();
 fill_2 FILLER_117_84 ();
 fill_1 FILLER_117_86 ();
 fill_1 FILLER_117_113 ();
 fill_2 FILLER_117_154 ();
 fill_4 FILLER_117_210 ();
 fill_1 FILLER_117_214 ();
 fill_2 FILLER_117_222 ();
 fill_4 FILLER_117_275 ();
 fill_1 FILLER_117_279 ();
 fill_1 FILLER_117_281 ();
 fill_2 FILLER_117_287 ();
 fill_1 FILLER_117_289 ();
 fill_4 FILLER_117_330 ();
 fill_2 FILLER_117_334 ();
 fill_2 FILLER_117_352 ();
 fill_1 FILLER_117_354 ();
 fill_2 FILLER_117_373 ();
 fill_1 FILLER_117_380 ();
 fill_1 FILLER_117_391 ();
 fill_2 FILLER_117_407 ();
 fill_8 FILLER_117_418 ();
 fill_1 FILLER_117_439 ();
 fill_2 FILLER_117_453 ();
 fill_2 FILLER_117_460 ();
 fill_1 FILLER_117_474 ();
 fill_2 FILLER_117_490 ();
 fill_1 FILLER_117_535 ();
 fill_2 FILLER_117_551 ();
 fill_4 FILLER_117_561 ();
 fill_2 FILLER_117_565 ();
 fill_2 FILLER_117_592 ();
 fill_2 FILLER_117_614 ();
 fill_2 FILLER_117_662 ();
 fill_1 FILLER_117_694 ();
 fill_1 FILLER_117_710 ();
 fill_1 FILLER_117_727 ();
 fill_1 FILLER_117_766 ();
 fill_2 FILLER_117_788 ();
 fill_1 FILLER_117_800 ();
 fill_4 FILLER_117_810 ();
 fill_2 FILLER_117_814 ();
 fill_2 FILLER_117_825 ();
 fill_2 FILLER_117_835 ();
 fill_2 FILLER_117_852 ();
 fill_1 FILLER_117_854 ();
 fill_1 FILLER_117_876 ();
 fill_1 FILLER_117_885 ();
 fill_2 FILLER_117_894 ();
 fill_8 FILLER_117_942 ();
 fill_2 FILLER_117_950 ();
 decap_12 FILLER_117_953 ();
 decap_12 FILLER_117_965 ();
 decap_12 FILLER_117_977 ();
 decap_12 FILLER_117_989 ();
 fill_4 FILLER_117_1001 ();
 fill_2 FILLER_117_1005 ();
 fill_1 FILLER_117_1007 ();
 decap_12 FILLER_117_1009 ();
 fill_4 FILLER_117_1021 ();
 fill_2 FILLER_117_1025 ();
 fill_1 FILLER_117_1027 ();
 decap_12 FILLER_118_3 ();
 decap_12 FILLER_118_15 ();
 fill_1 FILLER_118_27 ();
 decap_12 FILLER_118_29 ();
 decap_12 FILLER_118_41 ();
 fill_8 FILLER_118_53 ();
 fill_1 FILLER_118_61 ();
 fill_2 FILLER_118_82 ();
 fill_2 FILLER_118_105 ();
 fill_1 FILLER_118_150 ();
 fill_2 FILLER_118_201 ();
 fill_4 FILLER_118_218 ();
 fill_4 FILLER_118_260 ();
 decap_12 FILLER_118_271 ();
 fill_8 FILLER_118_283 ();
 fill_1 FILLER_118_291 ();
 fill_2 FILLER_118_306 ();
 fill_2 FILLER_118_309 ();
 fill_4 FILLER_118_325 ();
 fill_2 FILLER_118_337 ();
 fill_2 FILLER_118_355 ();
 fill_1 FILLER_118_357 ();
 fill_1 FILLER_118_365 ();
 decap_12 FILLER_118_387 ();
 fill_1 FILLER_118_399 ();
 fill_4 FILLER_118_405 ();
 fill_1 FILLER_118_419 ();
 fill_2 FILLER_118_428 ();
 fill_2 FILLER_118_446 ();
 fill_2 FILLER_118_454 ();
 fill_1 FILLER_118_475 ();
 fill_2 FILLER_118_492 ();
 fill_1 FILLER_118_494 ();
 fill_4 FILLER_118_528 ();
 fill_4 FILLER_118_533 ();
 fill_4 FILLER_118_545 ();
 fill_2 FILLER_118_549 ();
 fill_2 FILLER_118_556 ();
 fill_1 FILLER_118_558 ();
 decap_12 FILLER_118_566 ();
 fill_1 FILLER_118_578 ();
 fill_4 FILLER_118_584 ();
 fill_1 FILLER_118_589 ();
 fill_2 FILLER_118_622 ();
 fill_2 FILLER_118_701 ();
 fill_2 FILLER_118_729 ();
 fill_1 FILLER_118_755 ();
 fill_1 FILLER_118_783 ();
 fill_1 FILLER_118_790 ();
 fill_2 FILLER_118_837 ();
 fill_1 FILLER_118_839 ();
 fill_4 FILLER_118_848 ();
 fill_1 FILLER_118_852 ();
 fill_1 FILLER_118_869 ();
 fill_2 FILLER_118_874 ();
 fill_4 FILLER_118_880 ();
 fill_1 FILLER_118_884 ();
 fill_4 FILLER_118_888 ();
 fill_8 FILLER_118_896 ();
 fill_8 FILLER_118_915 ();
 fill_1 FILLER_118_923 ();
 decap_12 FILLER_118_932 ();
 decap_12 FILLER_118_944 ();
 decap_12 FILLER_118_956 ();
 decap_12 FILLER_118_968 ();
 decap_12 FILLER_118_981 ();
 decap_12 FILLER_118_993 ();
 decap_12 FILLER_118_1005 ();
 decap_12 FILLER_118_1017 ();
 fill_4 FILLER_118_1029 ();
 fill_2 FILLER_118_1033 ();
 fill_1 FILLER_118_1035 ();
 fill_1 FILLER_118_1037 ();
 decap_12 FILLER_119_3 ();
 decap_12 FILLER_119_15 ();
 decap_12 FILLER_119_27 ();
 decap_12 FILLER_119_39 ();
 fill_4 FILLER_119_51 ();
 fill_1 FILLER_119_55 ();
 fill_2 FILLER_119_77 ();
 fill_1 FILLER_119_88 ();
 fill_2 FILLER_119_109 ();
 fill_1 FILLER_119_111 ();
 fill_2 FILLER_119_117 ();
 fill_4 FILLER_119_169 ();
 fill_2 FILLER_119_173 ();
 fill_1 FILLER_119_204 ();
 fill_2 FILLER_119_222 ();
 fill_1 FILLER_119_225 ();
 fill_1 FILLER_119_233 ();
 fill_4 FILLER_119_254 ();
 fill_2 FILLER_119_258 ();
 fill_1 FILLER_119_260 ();
 decap_12 FILLER_119_291 ();
 fill_2 FILLER_119_303 ();
 fill_1 FILLER_119_305 ();
 fill_4 FILLER_119_330 ();
 fill_2 FILLER_119_334 ();
 fill_2 FILLER_119_337 ();
 fill_1 FILLER_119_355 ();
 fill_8 FILLER_119_372 ();
 fill_2 FILLER_119_380 ();
 fill_1 FILLER_119_391 ();
 fill_2 FILLER_119_428 ();
 fill_1 FILLER_119_435 ();
 fill_1 FILLER_119_457 ();
 fill_1 FILLER_119_479 ();
 fill_2 FILLER_119_497 ();
 fill_2 FILLER_119_531 ();
 fill_2 FILLER_119_540 ();
 fill_1 FILLER_119_542 ();
 fill_1 FILLER_119_559 ();
 fill_1 FILLER_119_569 ();
 fill_1 FILLER_119_583 ();
 fill_1 FILLER_119_637 ();
 fill_1 FILLER_119_682 ();
 fill_2 FILLER_119_688 ();
 fill_1 FILLER_119_719 ();
 fill_1 FILLER_119_727 ();
 fill_2 FILLER_119_738 ();
 fill_1 FILLER_119_740 ();
 fill_4 FILLER_119_766 ();
 fill_2 FILLER_119_770 ();
 fill_2 FILLER_119_785 ();
 fill_2 FILLER_119_810 ();
 fill_1 FILLER_119_812 ();
 fill_2 FILLER_119_821 ();
 fill_1 FILLER_119_823 ();
 fill_1 FILLER_119_828 ();
 fill_4 FILLER_119_836 ();
 fill_8 FILLER_119_866 ();
 fill_1 FILLER_119_895 ();
 fill_4 FILLER_119_897 ();
 fill_4 FILLER_119_908 ();
 fill_2 FILLER_119_912 ();
 fill_1 FILLER_119_914 ();
 fill_8 FILLER_119_943 ();
 fill_1 FILLER_119_951 ();
 decap_12 FILLER_119_953 ();
 decap_12 FILLER_119_965 ();
 decap_12 FILLER_119_977 ();
 decap_12 FILLER_119_989 ();
 fill_4 FILLER_119_1001 ();
 fill_2 FILLER_119_1005 ();
 fill_1 FILLER_119_1007 ();
 decap_12 FILLER_119_1009 ();
 decap_12 FILLER_119_1021 ();
 fill_4 FILLER_119_1033 ();
 fill_1 FILLER_119_1037 ();
 decap_12 FILLER_120_3 ();
 decap_12 FILLER_120_15 ();
 fill_1 FILLER_120_27 ();
 decap_12 FILLER_120_29 ();
 fill_2 FILLER_120_41 ();
 fill_1 FILLER_120_43 ();
 fill_1 FILLER_120_73 ();
 fill_2 FILLER_120_82 ();
 fill_1 FILLER_120_146 ();
 fill_2 FILLER_120_160 ();
 fill_1 FILLER_120_162 ();
 fill_1 FILLER_120_179 ();
 fill_2 FILLER_120_197 ();
 fill_1 FILLER_120_266 ();
 fill_4 FILLER_120_302 ();
 fill_2 FILLER_120_306 ();
 fill_8 FILLER_120_309 ();
 fill_2 FILLER_120_317 ();
 fill_1 FILLER_120_319 ();
 fill_1 FILLER_120_336 ();
 fill_1 FILLER_120_350 ();
 fill_2 FILLER_120_372 ();
 fill_4 FILLER_120_377 ();
 decap_12 FILLER_120_394 ();
 fill_4 FILLER_120_406 ();
 fill_1 FILLER_120_410 ();
 fill_2 FILLER_120_414 ();
 fill_1 FILLER_120_416 ();
 fill_1 FILLER_120_421 ();
 fill_2 FILLER_120_446 ();
 fill_1 FILLER_120_477 ();
 fill_1 FILLER_120_486 ();
 fill_1 FILLER_120_494 ();
 fill_1 FILLER_120_522 ();
 fill_1 FILLER_120_531 ();
 fill_2 FILLER_120_553 ();
 fill_1 FILLER_120_574 ();
 fill_1 FILLER_120_582 ();
 fill_2 FILLER_120_589 ();
 fill_2 FILLER_120_600 ();
 fill_1 FILLER_120_633 ();
 fill_1 FILLER_120_643 ();
 fill_2 FILLER_120_698 ();
 fill_1 FILLER_120_701 ();
 fill_4 FILLER_120_715 ();
 fill_4 FILLER_120_735 ();
 fill_2 FILLER_120_739 ();
 fill_4 FILLER_120_750 ();
 fill_2 FILLER_120_754 ();
 fill_1 FILLER_120_757 ();
 fill_1 FILLER_120_773 ();
 fill_1 FILLER_120_785 ();
 fill_2 FILLER_120_791 ();
 fill_2 FILLER_120_809 ();
 fill_1 FILLER_120_811 ();
 fill_1 FILLER_120_813 ();
 fill_1 FILLER_120_817 ();
 fill_2 FILLER_120_827 ();
 fill_1 FILLER_120_829 ();
 fill_8 FILLER_120_857 ();
 fill_2 FILLER_120_865 ();
 fill_1 FILLER_120_867 ();
 fill_4 FILLER_120_869 ();
 fill_1 FILLER_120_873 ();
 fill_8 FILLER_120_879 ();
 fill_2 FILLER_120_887 ();
 fill_2 FILLER_120_896 ();
 fill_1 FILLER_120_898 ();
 decap_12 FILLER_120_904 ();
 fill_4 FILLER_120_916 ();
 fill_1 FILLER_120_920 ();
 decap_12 FILLER_120_946 ();
 decap_12 FILLER_120_958 ();
 fill_8 FILLER_120_970 ();
 fill_2 FILLER_120_978 ();
 decap_12 FILLER_120_981 ();
 decap_12 FILLER_120_993 ();
 decap_12 FILLER_120_1005 ();
 decap_12 FILLER_120_1017 ();
 fill_4 FILLER_120_1029 ();
 fill_2 FILLER_120_1033 ();
 fill_1 FILLER_120_1035 ();
 fill_1 FILLER_120_1037 ();
 decap_12 FILLER_121_3 ();
 decap_12 FILLER_121_15 ();
 decap_12 FILLER_121_27 ();
 fill_8 FILLER_121_48 ();
 fill_2 FILLER_121_57 ();
 fill_4 FILLER_121_86 ();
 fill_1 FILLER_121_90 ();
 fill_1 FILLER_121_111 ();
 fill_2 FILLER_121_153 ();
 fill_1 FILLER_121_167 ();
 fill_1 FILLER_121_176 ();
 fill_2 FILLER_121_197 ();
 fill_2 FILLER_121_206 ();
 fill_2 FILLER_121_221 ();
 fill_1 FILLER_121_223 ();
 fill_2 FILLER_121_248 ();
 fill_2 FILLER_121_271 ();
 fill_1 FILLER_121_279 ();
 fill_1 FILLER_121_285 ();
 fill_4 FILLER_121_317 ();
 fill_4 FILLER_121_332 ();
 fill_1 FILLER_121_344 ();
 fill_1 FILLER_121_354 ();
 fill_1 FILLER_121_360 ();
 fill_1 FILLER_121_368 ();
 fill_8 FILLER_121_375 ();
 fill_2 FILLER_121_383 ();
 fill_2 FILLER_121_400 ();
 fill_4 FILLER_121_405 ();
 fill_2 FILLER_121_409 ();
 fill_2 FILLER_121_434 ();
 fill_1 FILLER_121_470 ();
 fill_1 FILLER_121_477 ();
 fill_1 FILLER_121_503 ();
 fill_1 FILLER_121_518 ();
 fill_2 FILLER_121_537 ();
 fill_4 FILLER_121_554 ();
 fill_2 FILLER_121_558 ();
 fill_1 FILLER_121_601 ();
 fill_1 FILLER_121_615 ();
 fill_1 FILLER_121_622 ();
 fill_1 FILLER_121_649 ();
 fill_2 FILLER_121_670 ();
 fill_4 FILLER_121_682 ();
 fill_2 FILLER_121_686 ();
 fill_1 FILLER_121_688 ();
 fill_2 FILLER_121_692 ();
 fill_1 FILLER_121_705 ();
 fill_2 FILLER_121_725 ();
 fill_1 FILLER_121_727 ();
 fill_1 FILLER_121_729 ();
 fill_4 FILLER_121_758 ();
 fill_2 FILLER_121_762 ();
 fill_1 FILLER_121_764 ();
 fill_1 FILLER_121_771 ();
 fill_1 FILLER_121_783 ();
 fill_1 FILLER_121_785 ();
 fill_8 FILLER_121_798 ();
 fill_1 FILLER_121_833 ();
 fill_4 FILLER_121_847 ();
 fill_1 FILLER_121_851 ();
 fill_2 FILLER_121_859 ();
 fill_2 FILLER_121_868 ();
 fill_4 FILLER_121_892 ();
 fill_1 FILLER_121_903 ();
 fill_2 FILLER_121_932 ();
 fill_8 FILLER_121_942 ();
 fill_2 FILLER_121_950 ();
 decap_12 FILLER_121_953 ();
 decap_12 FILLER_121_965 ();
 decap_12 FILLER_121_977 ();
 decap_12 FILLER_121_989 ();
 fill_4 FILLER_121_1001 ();
 fill_2 FILLER_121_1005 ();
 fill_1 FILLER_121_1007 ();
 decap_12 FILLER_121_1009 ();
 decap_12 FILLER_121_1021 ();
 fill_4 FILLER_121_1033 ();
 fill_1 FILLER_121_1037 ();
 decap_12 FILLER_122_3 ();
 decap_12 FILLER_122_15 ();
 fill_1 FILLER_122_27 ();
 fill_4 FILLER_122_29 ();
 fill_1 FILLER_122_33 ();
 fill_4 FILLER_122_54 ();
 fill_1 FILLER_122_77 ();
 fill_4 FILLER_122_114 ();
 fill_1 FILLER_122_118 ();
 fill_2 FILLER_122_128 ();
 fill_1 FILLER_122_130 ();
 fill_2 FILLER_122_180 ();
 fill_1 FILLER_122_195 ();
 fill_2 FILLER_122_197 ();
 fill_1 FILLER_122_199 ();
 fill_1 FILLER_122_209 ();
 fill_1 FILLER_122_245 ();
 fill_2 FILLER_122_317 ();
 fill_1 FILLER_122_348 ();
 decap_12 FILLER_122_380 ();
 fill_8 FILLER_122_392 ();
 fill_1 FILLER_122_400 ();
 fill_2 FILLER_122_417 ();
 fill_1 FILLER_122_419 ();
 fill_4 FILLER_122_428 ();
 fill_2 FILLER_122_432 ();
 fill_1 FILLER_122_454 ();
 fill_2 FILLER_122_477 ();
 fill_2 FILLER_122_513 ();
 fill_2 FILLER_122_597 ();
 fill_1 FILLER_122_633 ();
 fill_1 FILLER_122_643 ();
 fill_4 FILLER_122_715 ();
 fill_1 FILLER_122_719 ();
 fill_8 FILLER_122_737 ();
 fill_1 FILLER_122_745 ();
 fill_1 FILLER_122_755 ();
 fill_2 FILLER_122_760 ();
 fill_2 FILLER_122_771 ();
 fill_1 FILLER_122_773 ();
 fill_8 FILLER_122_800 ();
 fill_1 FILLER_122_808 ();
 fill_1 FILLER_122_813 ();
 fill_2 FILLER_122_817 ();
 fill_1 FILLER_122_825 ();
 fill_8 FILLER_122_857 ();
 fill_2 FILLER_122_865 ();
 fill_1 FILLER_122_867 ();
 fill_8 FILLER_122_881 ();
 fill_1 FILLER_122_889 ();
 fill_2 FILLER_122_896 ();
 fill_4 FILLER_122_918 ();
 fill_2 FILLER_122_922 ();
 decap_12 FILLER_122_934 ();
 decap_12 FILLER_122_946 ();
 decap_12 FILLER_122_958 ();
 fill_8 FILLER_122_970 ();
 fill_2 FILLER_122_978 ();
 decap_12 FILLER_122_981 ();
 decap_12 FILLER_122_993 ();
 decap_12 FILLER_122_1005 ();
 decap_12 FILLER_122_1017 ();
 fill_4 FILLER_122_1029 ();
 fill_2 FILLER_122_1033 ();
 fill_1 FILLER_122_1035 ();
 fill_1 FILLER_122_1037 ();
 decap_12 FILLER_123_3 ();
 decap_12 FILLER_123_15 ();
 fill_2 FILLER_123_53 ();
 fill_1 FILLER_123_55 ();
 fill_1 FILLER_123_91 ();
 fill_1 FILLER_123_134 ();
 fill_4 FILLER_123_217 ();
 fill_2 FILLER_123_221 ();
 fill_1 FILLER_123_223 ();
 fill_1 FILLER_123_260 ();
 fill_2 FILLER_123_278 ();
 fill_2 FILLER_123_300 ();
 fill_2 FILLER_123_324 ();
 fill_4 FILLER_123_330 ();
 fill_2 FILLER_123_334 ();
 fill_2 FILLER_123_337 ();
 decap_12 FILLER_123_347 ();
 decap_12 FILLER_123_359 ();
 fill_4 FILLER_123_385 ();
 fill_2 FILLER_123_389 ();
 fill_1 FILLER_123_391 ();
 fill_4 FILLER_123_400 ();
 fill_2 FILLER_123_404 ();
 fill_1 FILLER_123_406 ();
 fill_4 FILLER_123_434 ();
 fill_2 FILLER_123_438 ();
 fill_1 FILLER_123_447 ();
 fill_2 FILLER_123_452 ();
 fill_2 FILLER_123_505 ();
 fill_8 FILLER_123_543 ();
 fill_1 FILLER_123_551 ();
 fill_1 FILLER_123_561 ();
 fill_2 FILLER_123_566 ();
 fill_1 FILLER_123_577 ();
 fill_2 FILLER_123_587 ();
 fill_1 FILLER_123_589 ();
 fill_1 FILLER_123_671 ();
 fill_1 FILLER_123_694 ();
 fill_2 FILLER_123_702 ();
 fill_1 FILLER_123_711 ();
 fill_2 FILLER_123_723 ();
 fill_2 FILLER_123_729 ();
 fill_1 FILLER_123_745 ();
 fill_1 FILLER_123_785 ();
 fill_2 FILLER_123_789 ();
 fill_2 FILLER_123_838 ();
 fill_2 FILLER_123_845 ();
 fill_8 FILLER_123_853 ();
 fill_2 FILLER_123_869 ();
 fill_1 FILLER_123_871 ();
 fill_1 FILLER_123_878 ();
 fill_2 FILLER_123_888 ();
 fill_8 FILLER_123_908 ();
 decap_12 FILLER_123_922 ();
 decap_12 FILLER_123_934 ();
 fill_4 FILLER_123_946 ();
 fill_2 FILLER_123_950 ();
 decap_12 FILLER_123_953 ();
 decap_12 FILLER_123_965 ();
 decap_12 FILLER_123_977 ();
 decap_12 FILLER_123_989 ();
 fill_4 FILLER_123_1001 ();
 fill_2 FILLER_123_1005 ();
 fill_1 FILLER_123_1007 ();
 decap_12 FILLER_123_1009 ();
 decap_12 FILLER_123_1021 ();
 fill_4 FILLER_123_1033 ();
 fill_1 FILLER_123_1037 ();
 decap_12 FILLER_124_3 ();
 decap_12 FILLER_124_15 ();
 fill_1 FILLER_124_27 ();
 fill_4 FILLER_124_29 ();
 fill_1 FILLER_124_33 ();
 fill_8 FILLER_124_43 ();
 fill_4 FILLER_124_80 ();
 fill_4 FILLER_124_92 ();
 fill_1 FILLER_124_96 ();
 fill_1 FILLER_124_139 ();
 fill_1 FILLER_124_169 ();
 fill_1 FILLER_124_195 ();
 fill_4 FILLER_124_224 ();
 fill_1 FILLER_124_228 ();
 fill_2 FILLER_124_253 ();
 fill_1 FILLER_124_272 ();
 fill_2 FILLER_124_293 ();
 fill_2 FILLER_124_298 ();
 fill_2 FILLER_124_306 ();
 fill_2 FILLER_124_317 ();
 fill_2 FILLER_124_326 ();
 fill_2 FILLER_124_355 ();
 fill_1 FILLER_124_357 ();
 fill_4 FILLER_124_365 ();
 fill_1 FILLER_124_369 ();
 fill_4 FILLER_124_373 ();
 fill_2 FILLER_124_377 ();
 fill_1 FILLER_124_379 ();
 decap_12 FILLER_124_385 ();
 fill_1 FILLER_124_397 ();
 fill_2 FILLER_124_409 ();
 fill_2 FILLER_124_418 ();
 fill_2 FILLER_124_421 ();
 fill_2 FILLER_124_477 ();
 fill_1 FILLER_124_537 ();
 fill_2 FILLER_124_577 ();
 fill_1 FILLER_124_587 ();
 fill_2 FILLER_124_607 ();
 fill_2 FILLER_124_682 ();
 fill_2 FILLER_124_692 ();
 fill_2 FILLER_124_701 ();
 fill_2 FILLER_124_710 ();
 fill_1 FILLER_124_722 ();
 fill_1 FILLER_124_730 ();
 fill_4 FILLER_124_738 ();
 fill_2 FILLER_124_742 ();
 fill_1 FILLER_124_744 ();
 fill_1 FILLER_124_755 ();
 fill_4 FILLER_124_757 ();
 decap_12 FILLER_124_768 ();
 fill_2 FILLER_124_780 ();
 fill_2 FILLER_124_810 ();
 fill_8 FILLER_124_840 ();
 fill_2 FILLER_124_848 ();
 fill_1 FILLER_124_850 ();
 fill_4 FILLER_124_863 ();
 fill_1 FILLER_124_867 ();
 fill_2 FILLER_124_872 ();
 fill_4 FILLER_124_884 ();
 fill_1 FILLER_124_888 ();
 fill_2 FILLER_124_899 ();
 fill_2 FILLER_124_915 ();
 fill_4 FILLER_124_932 ();
 fill_2 FILLER_124_936 ();
 fill_1 FILLER_124_938 ();
 decap_12 FILLER_124_944 ();
 fill_4 FILLER_124_956 ();
 fill_8 FILLER_124_969 ();
 fill_2 FILLER_124_977 ();
 fill_1 FILLER_124_979 ();
 decap_12 FILLER_124_981 ();
 decap_12 FILLER_124_993 ();
 decap_12 FILLER_124_1005 ();
 decap_12 FILLER_124_1017 ();
 fill_4 FILLER_124_1029 ();
 fill_2 FILLER_124_1033 ();
 fill_1 FILLER_124_1035 ();
 fill_1 FILLER_124_1037 ();
 decap_12 FILLER_125_3 ();
 fill_1 FILLER_125_15 ();
 fill_2 FILLER_125_57 ();
 fill_1 FILLER_125_59 ();
 fill_1 FILLER_125_67 ();
 fill_1 FILLER_125_88 ();
 fill_2 FILLER_125_113 ();
 fill_4 FILLER_125_135 ();
 fill_1 FILLER_125_139 ();
 fill_4 FILLER_125_149 ();
 fill_1 FILLER_125_153 ();
 fill_1 FILLER_125_169 ();
 fill_1 FILLER_125_223 ();
 fill_1 FILLER_125_253 ();
 fill_1 FILLER_125_279 ();
 fill_1 FILLER_125_297 ();
 fill_2 FILLER_125_333 ();
 fill_1 FILLER_125_335 ();
 fill_2 FILLER_125_361 ();
 fill_2 FILLER_125_375 ();
 fill_2 FILLER_125_390 ();
 decap_12 FILLER_125_393 ();
 fill_2 FILLER_125_405 ();
 fill_1 FILLER_125_407 ();
 fill_2 FILLER_125_417 ();
 fill_1 FILLER_125_419 ();
 fill_4 FILLER_125_427 ();
 fill_1 FILLER_125_444 ();
 fill_2 FILLER_125_449 ();
 fill_1 FILLER_125_482 ();
 fill_1 FILLER_125_503 ();
 fill_1 FILLER_125_505 ();
 fill_1 FILLER_125_510 ();
 fill_2 FILLER_125_550 ();
 fill_2 FILLER_125_614 ();
 fill_2 FILLER_125_657 ();
 fill_2 FILLER_125_681 ();
 fill_2 FILLER_125_693 ();
 fill_4 FILLER_125_704 ();
 fill_2 FILLER_125_708 ();
 fill_1 FILLER_125_727 ();
 fill_2 FILLER_125_736 ();
 fill_1 FILLER_125_748 ();
 fill_1 FILLER_125_764 ();
 fill_2 FILLER_125_838 ();
 fill_1 FILLER_125_855 ();
 fill_1 FILLER_125_868 ();
 fill_1 FILLER_125_895 ();
 decap_12 FILLER_125_901 ();
 decap_12 FILLER_125_913 ();
 fill_2 FILLER_125_925 ();
 decap_12 FILLER_125_975 ();
 decap_12 FILLER_125_987 ();
 fill_8 FILLER_125_999 ();
 fill_1 FILLER_125_1007 ();
 decap_12 FILLER_125_1009 ();
 decap_12 FILLER_125_1021 ();
 fill_4 FILLER_125_1033 ();
 fill_1 FILLER_125_1037 ();
 decap_12 FILLER_126_3 ();
 decap_12 FILLER_126_15 ();
 fill_1 FILLER_126_27 ();
 fill_2 FILLER_126_29 ();
 fill_1 FILLER_126_31 ();
 fill_2 FILLER_126_41 ();
 fill_2 FILLER_126_137 ();
 fill_1 FILLER_126_139 ();
 fill_1 FILLER_126_150 ();
 fill_1 FILLER_126_195 ();
 fill_1 FILLER_126_197 ();
 fill_1 FILLER_126_217 ();
 fill_1 FILLER_126_309 ();
 fill_1 FILLER_126_339 ();
 fill_1 FILLER_126_368 ();
 fill_1 FILLER_126_378 ();
 fill_2 FILLER_126_417 ();
 fill_1 FILLER_126_419 ();
 fill_2 FILLER_126_437 ();
 fill_2 FILLER_126_465 ();
 fill_1 FILLER_126_486 ();
 fill_2 FILLER_126_499 ();
 fill_2 FILLER_126_533 ();
 fill_1 FILLER_126_593 ();
 fill_1 FILLER_126_621 ();
 fill_1 FILLER_126_721 ();
 fill_1 FILLER_126_742 ();
 fill_4 FILLER_126_750 ();
 fill_2 FILLER_126_754 ();
 fill_2 FILLER_126_799 ();
 fill_1 FILLER_126_811 ();
 fill_2 FILLER_126_845 ();
 fill_2 FILLER_126_850 ();
 fill_2 FILLER_126_866 ();
 fill_1 FILLER_126_874 ();
 fill_8 FILLER_126_878 ();
 fill_2 FILLER_126_886 ();
 fill_4 FILLER_126_898 ();
 fill_1 FILLER_126_902 ();
 fill_4 FILLER_126_910 ();
 fill_2 FILLER_126_921 ();
 fill_1 FILLER_126_923 ();
 fill_4 FILLER_126_925 ();
 fill_2 FILLER_126_945 ();
 fill_8 FILLER_126_951 ();
 fill_2 FILLER_126_959 ();
 fill_1 FILLER_126_961 ();
 fill_8 FILLER_126_971 ();
 fill_1 FILLER_126_979 ();
 decap_12 FILLER_126_981 ();
 decap_12 FILLER_126_993 ();
 decap_12 FILLER_126_1005 ();
 decap_12 FILLER_126_1017 ();
 fill_2 FILLER_126_1029 ();
 fill_1 FILLER_126_1031 ();
 fill_1 FILLER_126_1037 ();
 decap_12 FILLER_127_3 ();
 fill_8 FILLER_127_15 ();
 fill_2 FILLER_127_23 ();
 fill_1 FILLER_127_25 ();
 fill_4 FILLER_127_52 ();
 fill_1 FILLER_127_57 ();
 fill_2 FILLER_127_67 ();
 fill_1 FILLER_127_69 ();
 fill_4 FILLER_127_85 ();
 fill_4 FILLER_127_169 ();
 fill_1 FILLER_127_225 ();
 fill_1 FILLER_127_235 ();
 fill_1 FILLER_127_316 ();
 fill_2 FILLER_127_340 ();
 fill_1 FILLER_127_342 ();
 fill_8 FILLER_127_352 ();
 fill_1 FILLER_127_360 ();
 fill_1 FILLER_127_393 ();
 fill_2 FILLER_127_404 ();
 fill_1 FILLER_127_406 ();
 fill_2 FILLER_127_415 ();
 fill_8 FILLER_127_440 ();
 fill_4 FILLER_127_455 ();
 fill_2 FILLER_127_459 ();
 fill_2 FILLER_127_516 ();
 fill_2 FILLER_127_526 ();
 fill_2 FILLER_127_614 ();
 fill_2 FILLER_127_661 ();
 fill_1 FILLER_127_671 ();
 fill_2 FILLER_127_710 ();
 fill_2 FILLER_127_725 ();
 fill_1 FILLER_127_727 ();
 fill_2 FILLER_127_743 ();
 fill_1 FILLER_127_745 ();
 fill_4 FILLER_127_753 ();
 fill_4 FILLER_127_769 ();
 fill_2 FILLER_127_773 ();
 fill_2 FILLER_127_778 ();
 fill_1 FILLER_127_780 ();
 fill_1 FILLER_127_813 ();
 fill_1 FILLER_127_826 ();
 fill_1 FILLER_127_841 ();
 fill_2 FILLER_127_879 ();
 fill_1 FILLER_127_881 ();
 fill_1 FILLER_127_885 ();
 fill_2 FILLER_127_894 ();
 fill_1 FILLER_127_902 ();
 fill_1 FILLER_127_917 ();
 fill_2 FILLER_127_941 ();
 fill_2 FILLER_127_950 ();
 fill_4 FILLER_127_975 ();
 decap_12 FILLER_127_984 ();
 decap_12 FILLER_127_996 ();
 decap_12 FILLER_127_1009 ();
 decap_12 FILLER_127_1021 ();
 fill_4 FILLER_127_1033 ();
 fill_1 FILLER_127_1037 ();
 decap_12 FILLER_128_3 ();
 decap_12 FILLER_128_15 ();
 fill_1 FILLER_128_27 ();
 fill_2 FILLER_128_29 ();
 fill_1 FILLER_128_31 ();
 fill_1 FILLER_128_41 ();
 fill_2 FILLER_128_62 ();
 fill_1 FILLER_128_85 ();
 fill_1 FILLER_128_129 ();
 fill_2 FILLER_128_249 ();
 fill_1 FILLER_128_251 ();
 fill_1 FILLER_128_307 ();
 fill_4 FILLER_128_347 ();
 fill_2 FILLER_128_373 ();
 fill_2 FILLER_128_392 ();
 fill_1 FILLER_128_402 ();
 fill_1 FILLER_128_419 ();
 fill_1 FILLER_128_421 ();
 fill_1 FILLER_128_438 ();
 fill_8 FILLER_128_462 ();
 fill_2 FILLER_128_470 ();
 fill_1 FILLER_128_505 ();
 fill_1 FILLER_128_531 ();
 fill_1 FILLER_128_643 ();
 fill_2 FILLER_128_698 ();
 fill_1 FILLER_128_706 ();
 fill_2 FILLER_128_726 ();
 fill_1 FILLER_128_744 ();
 fill_2 FILLER_128_753 ();
 fill_1 FILLER_128_755 ();
 fill_1 FILLER_128_762 ();
 fill_2 FILLER_128_769 ();
 fill_2 FILLER_128_804 ();
 fill_1 FILLER_128_853 ();
 fill_1 FILLER_128_859 ();
 fill_2 FILLER_128_866 ();
 fill_4 FILLER_128_879 ();
 fill_2 FILLER_128_883 ();
 fill_1 FILLER_128_885 ();
 fill_4 FILLER_128_889 ();
 fill_8 FILLER_128_901 ();
 fill_1 FILLER_128_909 ();
 fill_2 FILLER_128_921 ();
 fill_1 FILLER_128_923 ();
 fill_4 FILLER_128_925 ();
 fill_1 FILLER_128_929 ();
 fill_4 FILLER_128_940 ();
 fill_2 FILLER_128_944 ();
 fill_4 FILLER_128_957 ();
 fill_2 FILLER_128_961 ();
 fill_1 FILLER_128_963 ();
 fill_2 FILLER_128_981 ();
 fill_1 FILLER_128_983 ();
 decap_12 FILLER_128_996 ();
 decap_12 FILLER_128_1008 ();
 decap_12 FILLER_128_1020 ();
 fill_4 FILLER_128_1032 ();
 fill_1 FILLER_128_1037 ();
 decap_12 FILLER_129_3 ();
 decap_12 FILLER_129_15 ();
 decap_12 FILLER_129_27 ();
 fill_4 FILLER_129_39 ();
 fill_1 FILLER_129_43 ();
 fill_4 FILLER_129_50 ();
 fill_2 FILLER_129_54 ();
 fill_2 FILLER_129_57 ();
 fill_1 FILLER_129_59 ();
 fill_2 FILLER_129_72 ();
 fill_1 FILLER_129_74 ();
 fill_4 FILLER_129_87 ();
 fill_1 FILLER_129_91 ();
 fill_2 FILLER_129_113 ();
 fill_2 FILLER_129_165 ();
 fill_1 FILLER_129_167 ();
 fill_1 FILLER_129_273 ();
 fill_1 FILLER_129_337 ();
 fill_1 FILLER_129_371 ();
 fill_1 FILLER_129_378 ();
 fill_2 FILLER_129_389 ();
 fill_1 FILLER_129_391 ();
 fill_1 FILLER_129_418 ();
 fill_2 FILLER_129_445 ();
 fill_1 FILLER_129_447 ();
 fill_1 FILLER_129_458 ();
 fill_4 FILLER_129_483 ();
 fill_2 FILLER_129_487 ();
 fill_1 FILLER_129_500 ();
 fill_1 FILLER_129_505 ();
 fill_2 FILLER_129_527 ();
 fill_2 FILLER_129_601 ();
 fill_1 FILLER_129_664 ();
 fill_1 FILLER_129_671 ();
 fill_1 FILLER_129_714 ();
 fill_1 FILLER_129_727 ();
 fill_1 FILLER_129_768 ();
 fill_2 FILLER_129_777 ();
 fill_1 FILLER_129_825 ();
 fill_2 FILLER_129_841 ();
 fill_1 FILLER_129_843 ();
 fill_1 FILLER_129_847 ();
 fill_4 FILLER_129_851 ();
 fill_1 FILLER_129_858 ();
 fill_4 FILLER_129_864 ();
 fill_2 FILLER_129_877 ();
 fill_4 FILLER_129_889 ();
 fill_2 FILLER_129_893 ();
 fill_1 FILLER_129_895 ();
 fill_4 FILLER_129_903 ();
 fill_1 FILLER_129_907 ();
 fill_2 FILLER_129_925 ();
 fill_8 FILLER_129_944 ();
 fill_2 FILLER_129_953 ();
 fill_8 FILLER_129_959 ();
 fill_1 FILLER_129_967 ();
 decap_12 FILLER_129_974 ();
 fill_2 FILLER_129_986 ();
 fill_1 FILLER_129_988 ();
 decap_12 FILLER_129_992 ();
 fill_4 FILLER_129_1004 ();
 decap_12 FILLER_129_1009 ();
 decap_12 FILLER_129_1021 ();
 fill_4 FILLER_129_1033 ();
 fill_1 FILLER_129_1037 ();
 decap_12 FILLER_130_3 ();
 decap_12 FILLER_130_15 ();
 fill_1 FILLER_130_27 ();
 fill_8 FILLER_130_29 ();
 fill_2 FILLER_130_66 ();
 fill_1 FILLER_130_83 ();
 fill_1 FILLER_130_106 ();
 fill_4 FILLER_130_148 ();
 fill_2 FILLER_130_194 ();
 fill_2 FILLER_130_203 ();
 fill_2 FILLER_130_231 ();
 fill_1 FILLER_130_233 ();
 fill_1 FILLER_130_243 ();
 fill_4 FILLER_130_253 ();
 fill_1 FILLER_130_266 ();
 fill_2 FILLER_130_309 ();
 fill_2 FILLER_130_348 ();
 fill_1 FILLER_130_350 ();
 fill_4 FILLER_130_381 ();
 fill_2 FILLER_130_385 ();
 decap_12 FILLER_130_421 ();
 fill_4 FILLER_130_433 ();
 fill_1 FILLER_130_437 ();
 fill_8 FILLER_130_448 ();
 fill_1 FILLER_130_456 ();
 fill_2 FILLER_130_471 ();
 fill_1 FILLER_130_477 ();
 fill_2 FILLER_130_484 ();
 fill_1 FILLER_130_528 ();
 fill_2 FILLER_130_533 ();
 fill_1 FILLER_130_567 ();
 fill_2 FILLER_130_597 ();
 fill_1 FILLER_130_599 ();
 fill_1 FILLER_130_643 ();
 fill_2 FILLER_130_687 ();
 fill_4 FILLER_130_728 ();
 fill_1 FILLER_130_732 ();
 fill_1 FILLER_130_739 ();
 fill_2 FILLER_130_747 ();
 fill_1 FILLER_130_755 ();
 fill_1 FILLER_130_769 ();
 decap_12 FILLER_130_773 ();
 fill_4 FILLER_130_785 ();
 fill_2 FILLER_130_789 ();
 fill_1 FILLER_130_791 ();
 fill_1 FILLER_130_850 ();
 fill_2 FILLER_130_869 ();
 fill_4 FILLER_130_883 ();
 fill_1 FILLER_130_887 ();
 fill_1 FILLER_130_909 ();
 fill_4 FILLER_130_918 ();
 fill_2 FILLER_130_922 ();
 fill_2 FILLER_130_925 ();
 fill_8 FILLER_130_935 ();
 fill_1 FILLER_130_943 ();
 fill_1 FILLER_130_947 ();
 fill_2 FILLER_130_955 ();
 fill_1 FILLER_130_957 ();
 fill_2 FILLER_130_970 ();
 fill_1 FILLER_130_989 ();
 decap_12 FILLER_130_1004 ();
 decap_12 FILLER_130_1016 ();
 fill_8 FILLER_130_1028 ();
 fill_1 FILLER_130_1037 ();
 decap_12 FILLER_131_3 ();
 decap_12 FILLER_131_15 ();
 fill_4 FILLER_131_27 ();
 fill_2 FILLER_131_31 ();
 fill_1 FILLER_131_33 ();
 fill_2 FILLER_131_54 ();
 fill_4 FILLER_131_57 ();
 fill_2 FILLER_131_89 ();
 fill_1 FILLER_131_104 ();
 fill_1 FILLER_131_138 ();
 fill_2 FILLER_131_178 ();
 fill_1 FILLER_131_196 ();
 fill_1 FILLER_131_217 ();
 fill_4 FILLER_131_225 ();
 fill_4 FILLER_131_249 ();
 fill_2 FILLER_131_269 ();
 fill_1 FILLER_131_302 ();
 fill_2 FILLER_131_334 ();
 fill_1 FILLER_131_375 ();
 decap_12 FILLER_131_407 ();
 fill_4 FILLER_131_419 ();
 decap_12 FILLER_131_430 ();
 fill_4 FILLER_131_442 ();
 fill_2 FILLER_131_446 ();
 fill_4 FILLER_131_455 ();
 fill_4 FILLER_131_467 ();
 fill_1 FILLER_131_471 ();
 decap_12 FILLER_131_475 ();
 decap_12 FILLER_131_487 ();
 fill_4 FILLER_131_499 ();
 fill_1 FILLER_131_503 ();
 fill_4 FILLER_131_513 ();
 fill_2 FILLER_131_523 ();
 fill_1 FILLER_131_528 ();
 fill_2 FILLER_131_536 ();
 fill_1 FILLER_131_559 ();
 fill_1 FILLER_131_655 ();
 fill_2 FILLER_131_673 ();
 fill_1 FILLER_131_691 ();
 fill_1 FILLER_131_729 ();
 fill_1 FILLER_131_737 ();
 fill_2 FILLER_131_745 ();
 fill_1 FILLER_131_747 ();
 fill_1 FILLER_131_783 ();
 fill_1 FILLER_131_848 ();
 fill_1 FILLER_131_856 ();
 fill_4 FILLER_131_860 ();
 fill_2 FILLER_131_864 ();
 fill_8 FILLER_131_869 ();
 decap_12 FILLER_131_883 ();
 fill_1 FILLER_131_895 ();
 fill_1 FILLER_131_904 ();
 fill_2 FILLER_131_916 ();
 fill_1 FILLER_131_918 ();
 fill_2 FILLER_131_933 ();
 fill_2 FILLER_131_949 ();
 fill_1 FILLER_131_951 ();
 fill_2 FILLER_131_953 ();
 fill_1 FILLER_131_955 ();
 fill_4 FILLER_131_960 ();
 fill_1 FILLER_131_964 ();
 fill_2 FILLER_131_978 ();
 fill_1 FILLER_131_1007 ();
 decap_12 FILLER_131_1009 ();
 decap_12 FILLER_131_1021 ();
 fill_4 FILLER_131_1033 ();
 fill_1 FILLER_131_1037 ();
 fill_4 FILLER_132_3 ();
 fill_1 FILLER_132_7 ();
 fill_8 FILLER_132_38 ();
 fill_4 FILLER_132_52 ();
 fill_2 FILLER_132_56 ();
 fill_4 FILLER_132_115 ();
 fill_1 FILLER_132_139 ();
 fill_1 FILLER_132_141 ();
 fill_2 FILLER_132_174 ();
 fill_4 FILLER_132_215 ();
 fill_1 FILLER_132_251 ();
 fill_2 FILLER_132_269 ();
 fill_1 FILLER_132_307 ();
 fill_1 FILLER_132_329 ();
 fill_2 FILLER_132_336 ();
 fill_2 FILLER_132_344 ();
 fill_1 FILLER_132_346 ();
 fill_1 FILLER_132_363 ();
 fill_2 FILLER_132_365 ();
 fill_8 FILLER_132_383 ();
 fill_2 FILLER_132_391 ();
 fill_1 FILLER_132_393 ();
 fill_2 FILLER_132_417 ();
 fill_1 FILLER_132_419 ();
 fill_8 FILLER_132_421 ();
 fill_2 FILLER_132_429 ();
 fill_1 FILLER_132_431 ();
 decap_12 FILLER_132_439 ();
 decap_12 FILLER_132_451 ();
 decap_12 FILLER_132_463 ();
 fill_1 FILLER_132_475 ();
 decap_12 FILLER_132_482 ();
 fill_4 FILLER_132_494 ();
 fill_8 FILLER_132_506 ();
 fill_4 FILLER_132_519 ();
 fill_2 FILLER_132_526 ();
 fill_1 FILLER_132_528 ();
 fill_2 FILLER_132_533 ();
 fill_1 FILLER_132_535 ();
 fill_1 FILLER_132_563 ();
 fill_1 FILLER_132_634 ();
 fill_1 FILLER_132_643 ();
 fill_1 FILLER_132_645 ();
 fill_1 FILLER_132_711 ();
 fill_4 FILLER_132_728 ();
 fill_8 FILLER_132_740 ();
 fill_4 FILLER_132_751 ();
 fill_1 FILLER_132_755 ();
 fill_2 FILLER_132_757 ();
 fill_4 FILLER_132_779 ();
 fill_2 FILLER_132_833 ();
 fill_4 FILLER_132_844 ();
 decap_12 FILLER_132_851 ();
 fill_4 FILLER_132_863 ();
 fill_1 FILLER_132_867 ();
 fill_1 FILLER_132_895 ();
 decap_12 FILLER_132_903 ();
 fill_8 FILLER_132_915 ();
 fill_1 FILLER_132_923 ();
 fill_8 FILLER_132_933 ();
 fill_4 FILLER_132_967 ();
 fill_2 FILLER_132_971 ();
 fill_1 FILLER_132_973 ();
 fill_1 FILLER_132_979 ();
 fill_2 FILLER_132_981 ();
 fill_1 FILLER_132_983 ();
 fill_2 FILLER_132_990 ();
 decap_12 FILLER_132_998 ();
 decap_12 FILLER_132_1010 ();
 decap_12 FILLER_132_1022 ();
 fill_2 FILLER_132_1034 ();
 fill_1 FILLER_132_1037 ();
 decap_12 FILLER_133_3 ();
 fill_1 FILLER_133_55 ();
 fill_2 FILLER_133_93 ();
 fill_1 FILLER_133_101 ();
 fill_2 FILLER_133_113 ();
 fill_1 FILLER_133_115 ();
 fill_2 FILLER_133_133 ();
 fill_1 FILLER_133_135 ();
 fill_2 FILLER_133_144 ();
 fill_1 FILLER_133_146 ();
 fill_1 FILLER_133_175 ();
 fill_2 FILLER_133_192 ();
 fill_1 FILLER_133_194 ();
 fill_2 FILLER_133_253 ();
 fill_1 FILLER_133_255 ();
 fill_2 FILLER_133_265 ();
 fill_1 FILLER_133_267 ();
 fill_4 FILLER_133_276 ();
 fill_4 FILLER_133_281 ();
 fill_4 FILLER_133_301 ();
 fill_1 FILLER_133_305 ();
 fill_1 FILLER_133_326 ();
 fill_1 FILLER_133_373 ();
 fill_2 FILLER_133_390 ();
 fill_8 FILLER_133_407 ();
 fill_2 FILLER_133_415 ();
 fill_1 FILLER_133_417 ();
 decap_12 FILLER_133_425 ();
 fill_4 FILLER_133_437 ();
 fill_2 FILLER_133_441 ();
 fill_4 FILLER_133_449 ();
 fill_2 FILLER_133_453 ();
 fill_1 FILLER_133_458 ();
 fill_2 FILLER_133_470 ();
 fill_1 FILLER_133_472 ();
 fill_8 FILLER_133_478 ();
 fill_1 FILLER_133_486 ();
 fill_2 FILLER_133_502 ();
 fill_8 FILLER_133_505 ();
 fill_4 FILLER_133_518 ();
 fill_2 FILLER_133_530 ();
 fill_1 FILLER_133_532 ();
 fill_2 FILLER_133_561 ();
 fill_1 FILLER_133_563 ();
 fill_1 FILLER_133_609 ();
 fill_1 FILLER_133_671 ();
 fill_1 FILLER_133_685 ();
 fill_1 FILLER_133_702 ();
 fill_2 FILLER_133_710 ();
 fill_1 FILLER_133_727 ();
 fill_1 FILLER_133_729 ();
 fill_2 FILLER_133_752 ();
 fill_1 FILLER_133_762 ();
 fill_4 FILLER_133_766 ();
 fill_2 FILLER_133_775 ();
 fill_1 FILLER_133_777 ();
 fill_2 FILLER_133_781 ();
 fill_1 FILLER_133_783 ();
 fill_2 FILLER_133_828 ();
 fill_2 FILLER_133_838 ();
 fill_2 FILLER_133_848 ();
 fill_1 FILLER_133_863 ();
 fill_2 FILLER_133_883 ();
 fill_1 FILLER_133_895 ();
 fill_1 FILLER_133_921 ();
 fill_1 FILLER_133_935 ();
 fill_2 FILLER_133_943 ();
 fill_1 FILLER_133_945 ();
 fill_2 FILLER_133_949 ();
 fill_1 FILLER_133_951 ();
 fill_1 FILLER_133_953 ();
 fill_4 FILLER_133_962 ();
 fill_2 FILLER_133_966 ();
 fill_1 FILLER_133_968 ();
 fill_4 FILLER_133_981 ();
 fill_2 FILLER_133_985 ();
 fill_1 FILLER_133_987 ();
 fill_4 FILLER_133_1003 ();
 fill_1 FILLER_133_1007 ();
 decap_12 FILLER_133_1009 ();
 decap_12 FILLER_133_1021 ();
 fill_4 FILLER_133_1033 ();
 fill_1 FILLER_133_1037 ();
 decap_12 FILLER_134_3 ();
 fill_4 FILLER_134_15 ();
 fill_1 FILLER_134_78 ();
 fill_2 FILLER_134_85 ();
 fill_1 FILLER_134_119 ();
 fill_1 FILLER_134_134 ();
 fill_2 FILLER_134_141 ();
 fill_4 FILLER_134_197 ();
 fill_2 FILLER_134_210 ();
 fill_1 FILLER_134_221 ();
 fill_2 FILLER_134_242 ();
 fill_2 FILLER_134_253 ();
 fill_4 FILLER_134_303 ();
 fill_1 FILLER_134_307 ();
 fill_8 FILLER_134_309 ();
 decap_12 FILLER_134_326 ();
 fill_1 FILLER_134_338 ();
 fill_2 FILLER_134_365 ();
 fill_1 FILLER_134_367 ();
 fill_4 FILLER_134_376 ();
 fill_8 FILLER_134_398 ();
 fill_1 FILLER_134_406 ();
 fill_8 FILLER_134_411 ();
 fill_1 FILLER_134_419 ();
 fill_8 FILLER_134_421 ();
 fill_2 FILLER_134_429 ();
 decap_12 FILLER_134_438 ();
 fill_4 FILLER_134_450 ();
 fill_2 FILLER_134_454 ();
 decap_12 FILLER_134_462 ();
 fill_2 FILLER_134_474 ();
 fill_4 FILLER_134_483 ();
 decap_12 FILLER_134_493 ();
 decap_12 FILLER_134_510 ();
 fill_8 FILLER_134_522 ();
 fill_2 FILLER_134_530 ();
 decap_12 FILLER_134_533 ();
 fill_2 FILLER_134_545 ();
 fill_1 FILLER_134_547 ();
 fill_2 FILLER_134_551 ();
 fill_1 FILLER_134_553 ();
 fill_8 FILLER_134_560 ();
 fill_1 FILLER_134_580 ();
 fill_2 FILLER_134_604 ();
 fill_1 FILLER_134_640 ();
 fill_1 FILLER_134_657 ();
 decap_12 FILLER_134_785 ();
 fill_2 FILLER_134_797 ();
 fill_2 FILLER_134_828 ();
 fill_1 FILLER_134_846 ();
 fill_4 FILLER_134_864 ();
 fill_4 FILLER_134_877 ();
 fill_1 FILLER_134_881 ();
 fill_4 FILLER_134_887 ();
 fill_1 FILLER_134_891 ();
 fill_2 FILLER_134_895 ();
 fill_1 FILLER_134_897 ();
 fill_8 FILLER_134_904 ();
 fill_2 FILLER_134_912 ();
 fill_1 FILLER_134_914 ();
 fill_2 FILLER_134_933 ();
 fill_1 FILLER_134_935 ();
 fill_4 FILLER_134_941 ();
 fill_1 FILLER_134_967 ();
 fill_4 FILLER_134_975 ();
 fill_1 FILLER_134_979 ();
 fill_1 FILLER_134_990 ();
 fill_1 FILLER_134_994 ();
 decap_12 FILLER_134_1010 ();
 decap_12 FILLER_134_1022 ();
 fill_2 FILLER_134_1034 ();
 fill_1 FILLER_134_1037 ();
 decap_12 FILLER_135_3 ();
 fill_4 FILLER_135_35 ();
 fill_2 FILLER_135_39 ();
 fill_1 FILLER_135_41 ();
 fill_4 FILLER_135_51 ();
 fill_1 FILLER_135_55 ();
 fill_2 FILLER_135_57 ();
 fill_4 FILLER_135_68 ();
 fill_1 FILLER_135_99 ();
 fill_1 FILLER_135_113 ();
 fill_2 FILLER_135_166 ();
 fill_1 FILLER_135_183 ();
 fill_2 FILLER_135_225 ();
 fill_2 FILLER_135_236 ();
 fill_2 FILLER_135_258 ();
 fill_1 FILLER_135_260 ();
 fill_1 FILLER_135_279 ();
 fill_2 FILLER_135_289 ();
 fill_1 FILLER_135_291 ();
 fill_4 FILLER_135_332 ();
 fill_2 FILLER_135_357 ();
 fill_2 FILLER_135_381 ();
 fill_1 FILLER_135_391 ();
 decap_12 FILLER_135_393 ();
 fill_8 FILLER_135_405 ();
 fill_2 FILLER_135_413 ();
 fill_8 FILLER_135_429 ();
 fill_2 FILLER_135_437 ();
 fill_1 FILLER_135_439 ();
 fill_2 FILLER_135_445 ();
 fill_1 FILLER_135_447 ();
 fill_1 FILLER_135_449 ();
 fill_1 FILLER_135_456 ();
 fill_2 FILLER_135_473 ();
 fill_1 FILLER_135_488 ();
 fill_2 FILLER_135_495 ();
 fill_1 FILLER_135_503 ();
 fill_8 FILLER_135_508 ();
 fill_2 FILLER_135_516 ();
 fill_4 FILLER_135_524 ();
 fill_2 FILLER_135_528 ();
 fill_1 FILLER_135_530 ();
 fill_4 FILLER_135_537 ();
 fill_1 FILLER_135_541 ();
 fill_8 FILLER_135_549 ();
 fill_2 FILLER_135_557 ();
 fill_1 FILLER_135_559 ();
 fill_8 FILLER_135_567 ();
 fill_2 FILLER_135_575 ();
 fill_2 FILLER_135_588 ();
 fill_1 FILLER_135_590 ();
 fill_1 FILLER_135_597 ();
 fill_8 FILLER_135_629 ();
 fill_1 FILLER_135_637 ();
 fill_2 FILLER_135_664 ();
 fill_1 FILLER_135_666 ();
 fill_1 FILLER_135_671 ();
 fill_4 FILLER_135_673 ();
 fill_1 FILLER_135_677 ();
 fill_2 FILLER_135_694 ();
 fill_2 FILLER_135_716 ();
 fill_1 FILLER_135_718 ();
 fill_2 FILLER_135_733 ();
 fill_1 FILLER_135_735 ();
 fill_4 FILLER_135_762 ();
 fill_2 FILLER_135_766 ();
 fill_4 FILLER_135_777 ();
 fill_2 FILLER_135_781 ();
 fill_1 FILLER_135_783 ();
 fill_2 FILLER_135_785 ();
 fill_1 FILLER_135_787 ();
 fill_2 FILLER_135_825 ();
 fill_1 FILLER_135_834 ();
 fill_1 FILLER_135_839 ();
 fill_2 FILLER_135_854 ();
 fill_1 FILLER_135_863 ();
 fill_4 FILLER_135_872 ();
 fill_2 FILLER_135_884 ();
 fill_4 FILLER_135_891 ();
 fill_1 FILLER_135_895 ();
 fill_4 FILLER_135_897 ();
 fill_2 FILLER_135_904 ();
 fill_8 FILLER_135_914 ();
 fill_4 FILLER_135_932 ();
 fill_2 FILLER_135_950 ();
 decap_12 FILLER_135_956 ();
 fill_4 FILLER_135_974 ();
 fill_2 FILLER_135_978 ();
 fill_1 FILLER_135_980 ();
 fill_8 FILLER_135_984 ();
 fill_2 FILLER_135_1005 ();
 fill_1 FILLER_135_1007 ();
 decap_12 FILLER_135_1009 ();
 decap_12 FILLER_135_1021 ();
 fill_1 FILLER_135_1033 ();
 decap_12 FILLER_136_3 ();
 decap_12 FILLER_136_15 ();
 fill_1 FILLER_136_27 ();
 fill_4 FILLER_136_29 ();
 fill_1 FILLER_136_33 ();
 fill_2 FILLER_136_63 ();
 fill_1 FILLER_136_65 ();
 fill_1 FILLER_136_78 ();
 fill_1 FILLER_136_89 ();
 fill_2 FILLER_136_137 ();
 fill_1 FILLER_136_139 ();
 fill_2 FILLER_136_141 ();
 fill_2 FILLER_136_152 ();
 fill_1 FILLER_136_174 ();
 fill_2 FILLER_136_182 ();
 fill_2 FILLER_136_206 ();
 fill_2 FILLER_136_217 ();
 fill_4 FILLER_136_224 ();
 fill_2 FILLER_136_228 ();
 fill_2 FILLER_136_238 ();
 fill_2 FILLER_136_249 ();
 fill_1 FILLER_136_251 ();
 fill_2 FILLER_136_253 ();
 fill_1 FILLER_136_255 ();
 fill_4 FILLER_136_287 ();
 fill_1 FILLER_136_291 ();
 fill_4 FILLER_136_309 ();
 fill_2 FILLER_136_313 ();
 fill_1 FILLER_136_315 ();
 fill_4 FILLER_136_334 ();
 fill_2 FILLER_136_338 ();
 fill_1 FILLER_136_340 ();
 fill_2 FILLER_136_365 ();
 fill_1 FILLER_136_380 ();
 fill_2 FILLER_136_402 ();
 fill_1 FILLER_136_404 ();
 fill_1 FILLER_136_408 ();
 fill_8 FILLER_136_412 ();
 fill_8 FILLER_136_421 ();
 fill_2 FILLER_136_429 ();
 fill_1 FILLER_136_431 ();
 decap_12 FILLER_136_441 ();
 fill_8 FILLER_136_453 ();
 fill_1 FILLER_136_461 ();
 fill_1 FILLER_136_475 ();
 fill_1 FILLER_136_490 ();
 fill_4 FILLER_136_495 ();
 fill_4 FILLER_136_503 ();
 fill_2 FILLER_136_507 ();
 fill_1 FILLER_136_509 ();
 fill_4 FILLER_136_528 ();
 decap_12 FILLER_136_533 ();
 fill_2 FILLER_136_545 ();
 fill_1 FILLER_136_547 ();
 fill_2 FILLER_136_571 ();
 fill_1 FILLER_136_573 ();
 fill_2 FILLER_136_586 ();
 fill_4 FILLER_136_589 ();
 fill_1 FILLER_136_603 ();
 fill_4 FILLER_136_630 ();
 fill_2 FILLER_136_634 ();
 fill_4 FILLER_136_640 ();
 decap_12 FILLER_136_645 ();
 decap_12 FILLER_136_657 ();
 decap_12 FILLER_136_669 ();
 fill_8 FILLER_136_681 ();
 fill_1 FILLER_136_689 ();
 fill_4 FILLER_136_693 ();
 fill_2 FILLER_136_697 ();
 fill_1 FILLER_136_699 ();
 fill_1 FILLER_136_704 ();
 fill_1 FILLER_136_709 ();
 fill_2 FILLER_136_730 ();
 fill_2 FILLER_136_749 ();
 fill_2 FILLER_136_766 ();
 fill_4 FILLER_136_802 ();
 fill_1 FILLER_136_813 ();
 fill_1 FILLER_136_838 ();
 fill_4 FILLER_136_846 ();
 fill_1 FILLER_136_850 ();
 fill_1 FILLER_136_859 ();
 fill_2 FILLER_136_866 ();
 fill_2 FILLER_136_869 ();
 fill_1 FILLER_136_871 ();
 fill_2 FILLER_136_879 ();
 fill_1 FILLER_136_881 ();
 fill_2 FILLER_136_895 ();
 fill_4 FILLER_136_900 ();
 fill_2 FILLER_136_904 ();
 fill_2 FILLER_136_916 ();
 fill_2 FILLER_136_925 ();
 fill_1 FILLER_136_927 ();
 fill_2 FILLER_136_933 ();
 fill_4 FILLER_136_941 ();
 fill_1 FILLER_136_945 ();
 fill_8 FILLER_136_954 ();
 fill_1 FILLER_136_962 ();
 decap_12 FILLER_136_996 ();
 decap_12 FILLER_136_1008 ();
 decap_12 FILLER_136_1020 ();
 fill_4 FILLER_136_1032 ();
 fill_1 FILLER_136_1037 ();
 fill_4 FILLER_137_57 ();
 fill_1 FILLER_137_85 ();
 fill_2 FILLER_137_98 ();
 fill_1 FILLER_137_113 ();
 fill_2 FILLER_137_155 ();
 fill_1 FILLER_137_182 ();
 fill_2 FILLER_137_197 ();
 fill_1 FILLER_137_199 ();
 fill_4 FILLER_137_220 ();
 fill_4 FILLER_137_225 ();
 fill_2 FILLER_137_229 ();
 fill_4 FILLER_137_260 ();
 fill_1 FILLER_137_271 ();
 fill_1 FILLER_137_279 ();
 fill_4 FILLER_137_281 ();
 fill_1 FILLER_137_285 ();
 fill_4 FILLER_137_302 ();
 fill_1 FILLER_137_306 ();
 fill_8 FILLER_137_337 ();
 fill_1 FILLER_137_354 ();
 fill_1 FILLER_137_391 ();
 decap_12 FILLER_137_393 ();
 decap_12 FILLER_137_405 ();
 fill_4 FILLER_137_417 ();
 decap_12 FILLER_137_424 ();
 decap_12 FILLER_137_436 ();
 decap_12 FILLER_137_458 ();
 fill_8 FILLER_137_470 ();
 fill_1 FILLER_137_478 ();
 fill_8 FILLER_137_494 ();
 fill_2 FILLER_137_502 ();
 fill_4 FILLER_137_511 ();
 fill_1 FILLER_137_515 ();
 fill_8 FILLER_137_525 ();
 fill_8 FILLER_137_551 ();
 fill_1 FILLER_137_559 ();
 fill_4 FILLER_137_561 ();
 fill_2 FILLER_137_565 ();
 fill_1 FILLER_137_567 ();
 fill_8 FILLER_137_574 ();
 fill_1 FILLER_137_588 ();
 fill_1 FILLER_137_597 ();
 decap_12 FILLER_137_631 ();
 fill_1 FILLER_137_643 ();
 fill_1 FILLER_137_662 ();
 fill_2 FILLER_137_673 ();
 fill_8 FILLER_137_682 ();
 fill_1 FILLER_137_690 ();
 fill_8 FILLER_137_729 ();
 fill_2 FILLER_137_737 ();
 fill_1 FILLER_137_739 ();
 fill_4 FILLER_137_779 ();
 fill_1 FILLER_137_783 ();
 fill_1 FILLER_137_813 ();
 fill_2 FILLER_137_841 ();
 fill_1 FILLER_137_843 ();
 fill_2 FILLER_137_852 ();
 fill_1 FILLER_137_854 ();
 fill_1 FILLER_137_867 ();
 fill_2 FILLER_137_885 ();
 fill_2 FILLER_137_894 ();
 fill_2 FILLER_137_972 ();
 fill_1 FILLER_137_974 ();
 fill_1 FILLER_137_986 ();
 fill_4 FILLER_137_992 ();
 fill_2 FILLER_137_996 ();
 fill_4 FILLER_137_1003 ();
 fill_1 FILLER_137_1007 ();
 decap_12 FILLER_137_1009 ();
 decap_12 FILLER_137_1021 ();
 fill_4 FILLER_137_1033 ();
 fill_1 FILLER_137_1037 ();
 decap_12 FILLER_138_3 ();
 fill_4 FILLER_138_15 ();
 fill_4 FILLER_138_29 ();
 fill_2 FILLER_138_82 ();
 fill_1 FILLER_138_132 ();
 fill_1 FILLER_138_184 ();
 fill_1 FILLER_138_206 ();
 fill_4 FILLER_138_247 ();
 fill_1 FILLER_138_251 ();
 fill_1 FILLER_138_259 ();
 fill_2 FILLER_138_269 ();
 fill_1 FILLER_138_271 ();
 fill_2 FILLER_138_286 ();
 fill_1 FILLER_138_307 ();
 fill_4 FILLER_138_309 ();
 fill_2 FILLER_138_322 ();
 fill_4 FILLER_138_344 ();
 fill_2 FILLER_138_348 ();
 fill_1 FILLER_138_350 ();
 fill_4 FILLER_138_374 ();
 fill_2 FILLER_138_378 ();
 fill_4 FILLER_138_396 ();
 fill_2 FILLER_138_400 ();
 fill_8 FILLER_138_409 ();
 fill_2 FILLER_138_417 ();
 fill_1 FILLER_138_419 ();
 fill_4 FILLER_138_424 ();
 decap_12 FILLER_138_443 ();
 fill_1 FILLER_138_455 ();
 fill_4 FILLER_138_501 ();
 fill_1 FILLER_138_505 ();
 decap_12 FILLER_138_519 ();
 fill_1 FILLER_138_531 ();
 fill_1 FILLER_138_533 ();
 fill_4 FILLER_138_539 ();
 fill_2 FILLER_138_543 ();
 fill_1 FILLER_138_568 ();
 fill_2 FILLER_138_585 ();
 fill_1 FILLER_138_587 ();
 fill_4 FILLER_138_597 ();
 fill_2 FILLER_138_601 ();
 fill_8 FILLER_138_619 ();
 fill_1 FILLER_138_627 ();
 fill_2 FILLER_138_633 ();
 fill_1 FILLER_138_635 ();
 fill_1 FILLER_138_643 ();
 fill_2 FILLER_138_653 ();
 decap_12 FILLER_138_664 ();
 fill_8 FILLER_138_676 ();
 fill_4 FILLER_138_687 ();
 fill_4 FILLER_138_694 ();
 fill_2 FILLER_138_698 ();
 fill_2 FILLER_138_704 ();
 fill_8 FILLER_138_747 ();
 fill_1 FILLER_138_755 ();
 fill_8 FILLER_138_757 ();
 fill_2 FILLER_138_765 ();
 fill_1 FILLER_138_767 ();
 fill_1 FILLER_138_811 ();
 fill_1 FILLER_138_857 ();
 fill_4 FILLER_138_864 ();
 fill_2 FILLER_138_869 ();
 fill_4 FILLER_138_908 ();
 fill_2 FILLER_138_912 ();
 fill_1 FILLER_138_914 ();
 fill_2 FILLER_138_922 ();
 fill_1 FILLER_138_932 ();
 fill_4 FILLER_138_941 ();
 fill_1 FILLER_138_945 ();
 fill_8 FILLER_138_953 ();
 fill_1 FILLER_138_961 ();
 fill_2 FILLER_138_969 ();
 fill_1 FILLER_138_979 ();
 fill_8 FILLER_138_981 ();
 fill_2 FILLER_138_989 ();
 fill_2 FILLER_138_994 ();
 decap_12 FILLER_138_999 ();
 decap_12 FILLER_138_1011 ();
 decap_12 FILLER_138_1023 ();
 fill_1 FILLER_138_1035 ();
 fill_1 FILLER_138_1037 ();
 fill_4 FILLER_139_3 ();
 fill_1 FILLER_139_7 ();
 fill_8 FILLER_139_48 ();
 fill_2 FILLER_139_57 ();
 fill_1 FILLER_139_59 ();
 fill_2 FILLER_139_100 ();
 fill_1 FILLER_139_111 ();
 fill_1 FILLER_139_113 ();
 fill_2 FILLER_139_159 ();
 fill_4 FILLER_139_169 ();
 fill_2 FILLER_139_173 ();
 fill_4 FILLER_139_184 ();
 fill_2 FILLER_139_188 ();
 fill_4 FILLER_139_210 ();
 fill_1 FILLER_139_214 ();
 fill_2 FILLER_139_278 ();
 fill_2 FILLER_139_281 ();
 fill_4 FILLER_139_310 ();
 fill_1 FILLER_139_314 ();
 fill_1 FILLER_139_335 ();
 fill_1 FILLER_139_357 ();
 fill_4 FILLER_139_385 ();
 fill_2 FILLER_139_389 ();
 fill_1 FILLER_139_391 ();
 fill_8 FILLER_139_396 ();
 decap_12 FILLER_139_411 ();
 decap_12 FILLER_139_423 ();
 fill_8 FILLER_139_435 ();
 fill_2 FILLER_139_443 ();
 fill_1 FILLER_139_456 ();
 fill_8 FILLER_139_470 ();
 fill_1 FILLER_139_478 ();
 fill_2 FILLER_139_482 ();
 fill_4 FILLER_139_498 ();
 fill_2 FILLER_139_502 ();
 fill_8 FILLER_139_505 ();
 fill_2 FILLER_139_513 ();
 fill_1 FILLER_139_515 ();
 fill_1 FILLER_139_520 ();
 fill_2 FILLER_139_527 ();
 fill_1 FILLER_139_529 ();
 decap_12 FILLER_139_533 ();
 fill_8 FILLER_139_545 ();
 fill_2 FILLER_139_553 ();
 fill_2 FILLER_139_558 ();
 fill_8 FILLER_139_561 ();
 fill_1 FILLER_139_569 ();
 fill_4 FILLER_139_578 ();
 fill_2 FILLER_139_582 ();
 fill_1 FILLER_139_584 ();
 fill_4 FILLER_139_598 ();
 fill_1 FILLER_139_602 ();
 fill_1 FILLER_139_607 ();
 fill_1 FILLER_139_615 ();
 fill_4 FILLER_139_628 ();
 fill_4 FILLER_139_638 ();
 fill_1 FILLER_139_642 ();
 fill_1 FILLER_139_650 ();
 fill_4 FILLER_139_665 ();
 fill_2 FILLER_139_669 ();
 fill_1 FILLER_139_671 ();
 fill_8 FILLER_139_676 ();
 fill_2 FILLER_139_697 ();
 fill_1 FILLER_139_699 ();
 fill_2 FILLER_139_778 ();
 fill_1 FILLER_139_780 ();
 fill_4 FILLER_139_855 ();
 fill_8 FILLER_139_864 ();
 fill_2 FILLER_139_872 ();
 fill_1 FILLER_139_874 ();
 fill_2 FILLER_139_897 ();
 fill_2 FILLER_139_906 ();
 fill_1 FILLER_139_908 ();
 fill_8 FILLER_139_912 ();
 fill_2 FILLER_139_920 ();
 fill_1 FILLER_139_922 ();
 fill_4 FILLER_139_930 ();
 fill_1 FILLER_139_939 ();
 fill_4 FILLER_139_945 ();
 fill_2 FILLER_139_949 ();
 fill_1 FILLER_139_951 ();
 fill_4 FILLER_139_953 ();
 fill_2 FILLER_139_957 ();
 fill_1 FILLER_139_959 ();
 fill_2 FILLER_139_971 ();
 fill_1 FILLER_139_973 ();
 fill_4 FILLER_139_1002 ();
 fill_2 FILLER_139_1006 ();
 decap_12 FILLER_139_1009 ();
 decap_12 FILLER_139_1021 ();
 fill_4 FILLER_139_1033 ();
 fill_1 FILLER_139_1037 ();
 decap_12 FILLER_140_3 ();
 decap_12 FILLER_140_15 ();
 fill_1 FILLER_140_27 ();
 fill_2 FILLER_140_29 ();
 fill_1 FILLER_140_31 ();
 fill_2 FILLER_140_61 ();
 fill_1 FILLER_140_63 ();
 fill_2 FILLER_140_85 ();
 fill_2 FILLER_140_137 ();
 fill_1 FILLER_140_139 ();
 fill_1 FILLER_140_154 ();
 fill_1 FILLER_140_229 ();
 fill_2 FILLER_140_250 ();
 fill_4 FILLER_140_253 ();
 fill_2 FILLER_140_257 ();
 fill_1 FILLER_140_259 ();
 fill_1 FILLER_140_292 ();
 fill_2 FILLER_140_306 ();
 fill_2 FILLER_140_338 ();
 fill_1 FILLER_140_365 ();
 fill_2 FILLER_140_380 ();
 decap_12 FILLER_140_407 ();
 fill_1 FILLER_140_419 ();
 fill_1 FILLER_140_421 ();
 fill_2 FILLER_140_425 ();
 fill_1 FILLER_140_427 ();
 fill_8 FILLER_140_431 ();
 fill_2 FILLER_140_439 ();
 fill_1 FILLER_140_446 ();
 fill_1 FILLER_140_454 ();
 fill_4 FILLER_140_460 ();
 fill_1 FILLER_140_464 ();
 fill_4 FILLER_140_484 ();
 fill_1 FILLER_140_488 ();
 fill_2 FILLER_140_497 ();
 fill_2 FILLER_140_510 ();
 fill_1 FILLER_140_516 ();
 fill_2 FILLER_140_523 ();
 fill_8 FILLER_140_550 ();
 fill_1 FILLER_140_558 ();
 fill_4 FILLER_140_582 ();
 fill_2 FILLER_140_586 ();
 fill_2 FILLER_140_589 ();
 fill_1 FILLER_140_591 ();
 fill_4 FILLER_140_622 ();
 fill_2 FILLER_140_626 ();
 fill_1 FILLER_140_628 ();
 fill_2 FILLER_140_642 ();
 fill_8 FILLER_140_645 ();
 fill_4 FILLER_140_675 ();
 fill_2 FILLER_140_679 ();
 fill_2 FILLER_140_697 ();
 fill_1 FILLER_140_699 ();
 fill_4 FILLER_140_725 ();
 fill_1 FILLER_140_729 ();
 fill_2 FILLER_140_735 ();
 fill_1 FILLER_140_746 ();
 fill_1 FILLER_140_813 ();
 fill_8 FILLER_140_851 ();
 fill_2 FILLER_140_859 ();
 fill_1 FILLER_140_861 ();
 fill_4 FILLER_140_901 ();
 fill_1 FILLER_140_905 ();
 fill_2 FILLER_140_909 ();
 fill_4 FILLER_140_919 ();
 fill_1 FILLER_140_923 ();
 fill_1 FILLER_140_941 ();
 fill_4 FILLER_140_957 ();
 fill_4 FILLER_140_970 ();
 fill_1 FILLER_140_974 ();
 fill_2 FILLER_140_991 ();
 fill_1 FILLER_140_993 ();
 decap_12 FILLER_140_1008 ();
 decap_12 FILLER_140_1020 ();
 fill_4 FILLER_140_1032 ();
 fill_1 FILLER_140_1037 ();
 decap_12 FILLER_141_3 ();
 decap_12 FILLER_141_15 ();
 fill_4 FILLER_141_27 ();
 fill_1 FILLER_141_31 ();
 fill_4 FILLER_141_52 ();
 fill_2 FILLER_141_66 ();
 fill_4 FILLER_141_117 ();
 fill_2 FILLER_141_121 ();
 fill_1 FILLER_141_129 ();
 fill_2 FILLER_141_150 ();
 fill_1 FILLER_141_169 ();
 fill_1 FILLER_141_190 ();
 fill_2 FILLER_141_211 ();
 fill_2 FILLER_141_216 ();
 fill_2 FILLER_141_234 ();
 fill_2 FILLER_141_290 ();
 fill_1 FILLER_141_292 ();
 fill_8 FILLER_141_302 ();
 fill_2 FILLER_141_330 ();
 fill_1 FILLER_141_332 ();
 fill_2 FILLER_141_373 ();
 fill_2 FILLER_141_407 ();
 fill_1 FILLER_141_409 ();
 fill_4 FILLER_141_416 ();
 fill_2 FILLER_141_420 ();
 fill_1 FILLER_141_422 ();
 fill_4 FILLER_141_433 ();
 fill_2 FILLER_141_437 ();
 fill_1 FILLER_141_439 ();
 fill_4 FILLER_141_443 ();
 fill_1 FILLER_141_447 ();
 fill_1 FILLER_141_449 ();
 fill_4 FILLER_141_463 ();
 fill_1 FILLER_141_473 ();
 decap_12 FILLER_141_480 ();
 fill_4 FILLER_141_492 ();
 fill_1 FILLER_141_496 ();
 fill_1 FILLER_141_503 ();
 decap_12 FILLER_141_514 ();
 fill_8 FILLER_141_526 ();
 fill_2 FILLER_141_541 ();
 fill_4 FILLER_141_547 ();
 fill_2 FILLER_141_551 ();
 fill_4 FILLER_141_556 ();
 fill_2 FILLER_141_561 ();
 fill_1 FILLER_141_583 ();
 fill_4 FILLER_141_588 ();
 fill_1 FILLER_141_592 ();
 fill_2 FILLER_141_597 ();
 decap_12 FILLER_141_602 ();
 fill_2 FILLER_141_614 ();
 fill_1 FILLER_141_617 ();
 fill_4 FILLER_141_630 ();
 fill_1 FILLER_141_642 ();
 fill_1 FILLER_141_651 ();
 fill_2 FILLER_141_660 ();
 fill_2 FILLER_141_670 ();
 fill_4 FILLER_141_689 ();
 fill_2 FILLER_141_693 ();
 fill_1 FILLER_141_695 ();
 fill_1 FILLER_141_727 ();
 fill_2 FILLER_141_782 ();
 fill_1 FILLER_141_802 ();
 fill_1 FILLER_141_839 ();
 fill_1 FILLER_141_864 ();
 fill_4 FILLER_141_872 ();
 fill_1 FILLER_141_876 ();
 fill_8 FILLER_141_888 ();
 fill_2 FILLER_141_900 ();
 fill_1 FILLER_141_902 ();
 fill_4 FILLER_141_918 ();
 fill_1 FILLER_141_922 ();
 fill_4 FILLER_141_930 ();
 fill_1 FILLER_141_934 ();
 fill_2 FILLER_141_938 ();
 fill_1 FILLER_141_940 ();
 fill_8 FILLER_141_944 ();
 fill_8 FILLER_141_964 ();
 fill_2 FILLER_141_972 ();
 fill_1 FILLER_141_974 ();
 fill_4 FILLER_141_979 ();
 fill_1 FILLER_141_983 ();
 fill_2 FILLER_141_993 ();
 fill_2 FILLER_141_1006 ();
 decap_12 FILLER_141_1009 ();
 decap_12 FILLER_141_1021 ();
 fill_4 FILLER_141_1033 ();
 fill_1 FILLER_141_1037 ();
 decap_12 FILLER_142_3 ();
 decap_12 FILLER_142_15 ();
 fill_1 FILLER_142_27 ();
 fill_2 FILLER_142_29 ();
 fill_1 FILLER_142_31 ();
 fill_2 FILLER_142_41 ();
 fill_1 FILLER_142_43 ();
 fill_2 FILLER_142_85 ();
 fill_1 FILLER_142_87 ();
 fill_4 FILLER_142_136 ();
 fill_4 FILLER_142_141 ();
 fill_1 FILLER_142_145 ();
 fill_1 FILLER_142_175 ();
 fill_1 FILLER_142_210 ();
 fill_2 FILLER_142_230 ();
 fill_1 FILLER_142_232 ();
 fill_1 FILLER_142_251 ();
 fill_1 FILLER_142_253 ();
 fill_4 FILLER_142_270 ();
 fill_2 FILLER_142_274 ();
 fill_1 FILLER_142_276 ();
 fill_2 FILLER_142_280 ();
 fill_1 FILLER_142_282 ();
 fill_2 FILLER_142_306 ();
 fill_2 FILLER_142_309 ();
 fill_1 FILLER_142_311 ();
 fill_4 FILLER_142_321 ();
 fill_1 FILLER_142_325 ();
 fill_2 FILLER_142_347 ();
 fill_8 FILLER_142_412 ();
 decap_12 FILLER_142_421 ();
 decap_12 FILLER_142_433 ();
 fill_4 FILLER_142_445 ();
 fill_2 FILLER_142_449 ();
 fill_4 FILLER_142_459 ();
 fill_2 FILLER_142_474 ();
 decap_12 FILLER_142_477 ();
 fill_2 FILLER_142_489 ();
 fill_2 FILLER_142_505 ();
 fill_1 FILLER_142_507 ();
 fill_2 FILLER_142_533 ();
 fill_1 FILLER_142_535 ();
 fill_2 FILLER_142_544 ();
 fill_2 FILLER_142_586 ();
 decap_12 FILLER_142_589 ();
 decap_12 FILLER_142_601 ();
 fill_2 FILLER_142_613 ();
 fill_1 FILLER_142_615 ();
 fill_4 FILLER_142_619 ();
 fill_2 FILLER_142_623 ();
 fill_1 FILLER_142_625 ();
 fill_4 FILLER_142_629 ();
 fill_1 FILLER_142_633 ();
 fill_4 FILLER_142_637 ();
 fill_2 FILLER_142_641 ();
 fill_1 FILLER_142_643 ();
 fill_2 FILLER_142_645 ();
 fill_1 FILLER_142_650 ();
 fill_4 FILLER_142_671 ();
 fill_2 FILLER_142_675 ();
 fill_1 FILLER_142_677 ();
 fill_2 FILLER_142_698 ();
 fill_2 FILLER_142_757 ();
 fill_1 FILLER_142_811 ();
 fill_2 FILLER_142_820 ();
 fill_4 FILLER_142_840 ();
 fill_2 FILLER_142_844 ();
 fill_2 FILLER_142_874 ();
 fill_4 FILLER_142_879 ();
 fill_1 FILLER_142_883 ();
 fill_1 FILLER_142_895 ();
 fill_8 FILLER_142_899 ();
 fill_2 FILLER_142_907 ();
 fill_2 FILLER_142_918 ();
 fill_1 FILLER_142_920 ();
 fill_1 FILLER_142_930 ();
 fill_2 FILLER_142_949 ();
 fill_1 FILLER_142_961 ();
 fill_4 FILLER_142_976 ();
 fill_8 FILLER_142_981 ();
 fill_2 FILLER_142_989 ();
 fill_1 FILLER_142_991 ();
 fill_8 FILLER_142_1002 ();
 decap_12 FILLER_142_1017 ();
 fill_4 FILLER_142_1029 ();
 fill_2 FILLER_142_1033 ();
 fill_1 FILLER_142_1035 ();
 fill_1 FILLER_142_1037 ();
 decap_12 FILLER_143_3 ();
 decap_12 FILLER_143_15 ();
 fill_8 FILLER_143_27 ();
 fill_2 FILLER_143_35 ();
 fill_1 FILLER_143_37 ();
 fill_4 FILLER_143_57 ();
 fill_4 FILLER_143_81 ();
 fill_2 FILLER_143_110 ();
 fill_4 FILLER_143_113 ();
 fill_2 FILLER_143_117 ();
 fill_4 FILLER_143_128 ();
 fill_1 FILLER_143_153 ();
 fill_2 FILLER_143_166 ();
 fill_1 FILLER_143_176 ();
 fill_2 FILLER_143_201 ();
 fill_1 FILLER_143_223 ();
 fill_1 FILLER_143_232 ();
 decap_12 FILLER_143_249 ();
 fill_2 FILLER_143_261 ();
 fill_1 FILLER_143_279 ();
 fill_2 FILLER_143_281 ();
 fill_4 FILLER_143_309 ();
 fill_1 FILLER_143_313 ();
 fill_4 FILLER_143_323 ();
 fill_2 FILLER_143_327 ();
 fill_2 FILLER_143_337 ();
 fill_2 FILLER_143_343 ();
 fill_2 FILLER_143_390 ();
 fill_4 FILLER_143_419 ();
 fill_1 FILLER_143_423 ();
 fill_2 FILLER_143_434 ();
 fill_8 FILLER_143_440 ();
 fill_2 FILLER_143_449 ();
 fill_1 FILLER_143_451 ();
 fill_1 FILLER_143_462 ();
 fill_2 FILLER_143_471 ();
 fill_1 FILLER_143_477 ();
 fill_4 FILLER_143_499 ();
 fill_1 FILLER_143_503 ();
 fill_8 FILLER_143_508 ();
 fill_1 FILLER_143_516 ();
 fill_2 FILLER_143_526 ();
 fill_2 FILLER_143_558 ();
 decap_12 FILLER_143_583 ();
 fill_2 FILLER_143_595 ();
 fill_2 FILLER_143_603 ();
 fill_1 FILLER_143_605 ();
 fill_2 FILLER_143_609 ();
 fill_1 FILLER_143_630 ();
 fill_1 FILLER_143_635 ();
 fill_2 FILLER_143_656 ();
 fill_8 FILLER_143_662 ();
 fill_2 FILLER_143_670 ();
 fill_1 FILLER_143_673 ();
 fill_4 FILLER_143_685 ();
 fill_2 FILLER_143_689 ();
 fill_4 FILLER_143_729 ();
 fill_1 FILLER_143_733 ();
 fill_2 FILLER_143_768 ();
 fill_1 FILLER_143_783 ();
 fill_1 FILLER_143_793 ();
 fill_4 FILLER_143_835 ();
 fill_1 FILLER_143_839 ();
 fill_2 FILLER_143_849 ();
 fill_1 FILLER_143_851 ();
 fill_2 FILLER_143_881 ();
 fill_1 FILLER_143_883 ();
 fill_8 FILLER_143_887 ();
 fill_1 FILLER_143_895 ();
 fill_8 FILLER_143_933 ();
 fill_1 FILLER_143_941 ();
 fill_1 FILLER_143_948 ();
 fill_1 FILLER_143_953 ();
 fill_2 FILLER_143_972 ();
 fill_1 FILLER_143_974 ();
 fill_1 FILLER_143_984 ();
 fill_4 FILLER_143_991 ();
 fill_2 FILLER_143_998 ();
 fill_4 FILLER_143_1034 ();
 decap_12 FILLER_144_3 ();
 decap_12 FILLER_144_15 ();
 fill_1 FILLER_144_27 ();
 fill_4 FILLER_144_29 ();
 fill_2 FILLER_144_33 ();
 fill_8 FILLER_144_76 ();
 fill_1 FILLER_144_105 ();
 fill_4 FILLER_144_135 ();
 fill_1 FILLER_144_139 ();
 fill_2 FILLER_144_161 ();
 fill_2 FILLER_144_197 ();
 fill_1 FILLER_144_221 ();
 fill_4 FILLER_144_263 ();
 fill_1 FILLER_144_267 ();
 fill_1 FILLER_144_272 ();
 fill_1 FILLER_144_296 ();
 fill_2 FILLER_144_306 ();
 fill_2 FILLER_144_309 ();
 fill_1 FILLER_144_363 ();
 fill_4 FILLER_144_387 ();
 fill_2 FILLER_144_391 ();
 fill_1 FILLER_144_419 ();
 fill_4 FILLER_144_424 ();
 fill_1 FILLER_144_428 ();
 fill_8 FILLER_144_432 ();
 fill_2 FILLER_144_440 ();
 fill_1 FILLER_144_442 ();
 decap_12 FILLER_144_454 ();
 fill_2 FILLER_144_466 ();
 fill_1 FILLER_144_468 ();
 decap_12 FILLER_144_477 ();
 fill_4 FILLER_144_489 ();
 fill_2 FILLER_144_493 ();
 fill_1 FILLER_144_495 ();
 fill_2 FILLER_144_512 ();
 fill_1 FILLER_144_514 ();
 fill_1 FILLER_144_522 ();
 fill_2 FILLER_144_530 ();
 fill_2 FILLER_144_533 ();
 fill_2 FILLER_144_566 ();
 fill_8 FILLER_144_579 ();
 fill_1 FILLER_144_587 ();
 fill_8 FILLER_144_597 ();
 fill_2 FILLER_144_605 ();
 fill_2 FILLER_144_631 ();
 fill_4 FILLER_144_645 ();
 fill_2 FILLER_144_649 ();
 fill_8 FILLER_144_657 ();
 fill_2 FILLER_144_665 ();
 fill_1 FILLER_144_667 ();
 fill_2 FILLER_144_697 ();
 fill_1 FILLER_144_699 ();
 fill_2 FILLER_144_710 ();
 fill_1 FILLER_144_755 ();
 fill_2 FILLER_144_768 ();
 fill_1 FILLER_144_783 ();
 fill_2 FILLER_144_801 ();
 fill_4 FILLER_144_862 ();
 fill_2 FILLER_144_866 ();
 fill_4 FILLER_144_876 ();
 fill_2 FILLER_144_880 ();
 fill_1 FILLER_144_882 ();
 fill_2 FILLER_144_889 ();
 fill_1 FILLER_144_891 ();
 fill_2 FILLER_144_907 ();
 fill_1 FILLER_144_923 ();
 fill_4 FILLER_144_932 ();
 fill_2 FILLER_144_936 ();
 fill_1 FILLER_144_938 ();
 fill_1 FILLER_144_949 ();
 fill_4 FILLER_144_956 ();
 fill_1 FILLER_144_960 ();
 fill_1 FILLER_144_970 ();
 fill_2 FILLER_144_978 ();
 fill_8 FILLER_144_981 ();
 fill_2 FILLER_144_989 ();
 fill_2 FILLER_144_1003 ();
 decap_12 FILLER_144_1015 ();
 fill_2 FILLER_144_1027 ();
 fill_1 FILLER_144_1029 ();
 fill_1 FILLER_144_1037 ();
 decap_12 FILLER_145_3 ();
 decap_12 FILLER_145_15 ();
 decap_12 FILLER_145_27 ();
 fill_4 FILLER_145_39 ();
 fill_1 FILLER_145_43 ();
 fill_2 FILLER_145_53 ();
 fill_1 FILLER_145_55 ();
 fill_2 FILLER_145_57 ();
 fill_1 FILLER_145_59 ();
 fill_2 FILLER_145_78 ();
 fill_1 FILLER_145_80 ();
 fill_2 FILLER_145_110 ();
 fill_4 FILLER_145_133 ();
 fill_2 FILLER_145_137 ();
 fill_4 FILLER_145_191 ();
 fill_1 FILLER_145_195 ();
 decap_12 FILLER_145_249 ();
 fill_2 FILLER_145_261 ();
 fill_1 FILLER_145_263 ();
 fill_4 FILLER_145_270 ();
 fill_2 FILLER_145_277 ();
 fill_1 FILLER_145_279 ();
 decap_12 FILLER_145_281 ();
 fill_8 FILLER_145_293 ();
 fill_2 FILLER_145_331 ();
 fill_4 FILLER_145_364 ();
 fill_2 FILLER_145_389 ();
 fill_1 FILLER_145_391 ();
 fill_1 FILLER_145_393 ();
 fill_1 FILLER_145_405 ();
 fill_1 FILLER_145_419 ();
 fill_1 FILLER_145_436 ();
 fill_2 FILLER_145_446 ();
 fill_4 FILLER_145_452 ();
 fill_2 FILLER_145_456 ();
 fill_8 FILLER_145_463 ();
 fill_2 FILLER_145_471 ();
 decap_12 FILLER_145_479 ();
 fill_8 FILLER_145_496 ();
 fill_2 FILLER_145_505 ();
 fill_1 FILLER_145_507 ();
 fill_2 FILLER_145_519 ();
 fill_1 FILLER_145_521 ();
 fill_2 FILLER_145_535 ();
 fill_1 FILLER_145_537 ();
 fill_4 FILLER_145_544 ();
 fill_1 FILLER_145_548 ();
 fill_2 FILLER_145_557 ();
 fill_1 FILLER_145_559 ();
 fill_2 FILLER_145_573 ();
 fill_1 FILLER_145_575 ();
 fill_2 FILLER_145_583 ();
 fill_1 FILLER_145_585 ();
 fill_8 FILLER_145_592 ();
 fill_2 FILLER_145_600 ();
 fill_4 FILLER_145_612 ();
 fill_4 FILLER_145_641 ();
 fill_1 FILLER_145_645 ();
 fill_1 FILLER_145_671 ();
 fill_4 FILLER_145_693 ();
 fill_1 FILLER_145_697 ();
 fill_2 FILLER_145_704 ();
 fill_2 FILLER_145_729 ();
 fill_2 FILLER_145_765 ();
 fill_1 FILLER_145_819 ();
 fill_2 FILLER_145_829 ();
 fill_1 FILLER_145_860 ();
 decap_12 FILLER_145_897 ();
 fill_2 FILLER_145_909 ();
 fill_4 FILLER_145_918 ();
 fill_8 FILLER_145_971 ();
 fill_2 FILLER_145_979 ();
 fill_1 FILLER_145_981 ();
 fill_2 FILLER_145_1006 ();
 decap_12 FILLER_145_1021 ();
 fill_4 FILLER_145_1033 ();
 fill_1 FILLER_145_1037 ();
 decap_12 FILLER_146_3 ();
 decap_12 FILLER_146_15 ();
 fill_1 FILLER_146_27 ();
 fill_8 FILLER_146_29 ();
 fill_1 FILLER_146_37 ();
 fill_2 FILLER_146_58 ();
 fill_1 FILLER_146_60 ();
 fill_2 FILLER_146_81 ();
 fill_1 FILLER_146_83 ();
 fill_2 FILLER_146_85 ();
 fill_1 FILLER_146_87 ();
 fill_2 FILLER_146_137 ();
 fill_1 FILLER_146_139 ();
 fill_4 FILLER_146_150 ();
 fill_2 FILLER_146_154 ();
 fill_1 FILLER_146_176 ();
 fill_2 FILLER_146_201 ();
 fill_8 FILLER_146_263 ();
 fill_2 FILLER_146_291 ();
 fill_1 FILLER_146_307 ();
 fill_2 FILLER_146_312 ();
 fill_1 FILLER_146_323 ();
 fill_2 FILLER_146_362 ();
 fill_2 FILLER_146_371 ();
 fill_1 FILLER_146_373 ();
 fill_2 FILLER_146_380 ();
 fill_1 FILLER_146_389 ();
 fill_4 FILLER_146_397 ();
 fill_2 FILLER_146_401 ();
 fill_4 FILLER_146_406 ();
 fill_2 FILLER_146_410 ();
 fill_4 FILLER_146_416 ();
 fill_4 FILLER_146_436 ();
 fill_2 FILLER_146_440 ();
 fill_1 FILLER_146_442 ();
 fill_4 FILLER_146_448 ();
 decap_12 FILLER_146_460 ();
 fill_4 FILLER_146_472 ();
 fill_2 FILLER_146_482 ();
 fill_1 FILLER_146_484 ();
 decap_12 FILLER_146_493 ();
 fill_4 FILLER_146_505 ();
 fill_4 FILLER_146_515 ();
 fill_2 FILLER_146_519 ();
 fill_2 FILLER_146_530 ();
 fill_2 FILLER_146_536 ();
 fill_2 FILLER_146_547 ();
 fill_1 FILLER_146_549 ();
 fill_2 FILLER_146_566 ();
 fill_2 FILLER_146_585 ();
 fill_1 FILLER_146_587 ();
 fill_1 FILLER_146_599 ();
 fill_2 FILLER_146_613 ();
 fill_1 FILLER_146_615 ();
 fill_4 FILLER_146_624 ();
 fill_2 FILLER_146_628 ();
 fill_1 FILLER_146_630 ();
 fill_1 FILLER_146_634 ();
 fill_2 FILLER_146_645 ();
 fill_2 FILLER_146_654 ();
 fill_1 FILLER_146_685 ();
 fill_4 FILLER_146_695 ();
 fill_1 FILLER_146_699 ();
 fill_1 FILLER_146_771 ();
 fill_2 FILLER_146_784 ();
 fill_1 FILLER_146_795 ();
 fill_1 FILLER_146_805 ();
 fill_1 FILLER_146_825 ();
 fill_2 FILLER_146_869 ();
 fill_2 FILLER_146_903 ();
 fill_4 FILLER_146_919 ();
 fill_1 FILLER_146_923 ();
 fill_1 FILLER_146_952 ();
 fill_2 FILLER_146_984 ();
 fill_1 FILLER_146_986 ();
 fill_2 FILLER_146_997 ();
 fill_1 FILLER_146_1008 ();
 fill_1 FILLER_146_1037 ();
 decap_12 FILLER_147_3 ();
 decap_12 FILLER_147_15 ();
 fill_8 FILLER_147_27 ();
 fill_2 FILLER_147_35 ();
 fill_1 FILLER_147_37 ();
 fill_4 FILLER_147_57 ();
 fill_4 FILLER_147_82 ();
 fill_2 FILLER_147_86 ();
 fill_4 FILLER_147_108 ();
 fill_2 FILLER_147_119 ();
 fill_1 FILLER_147_130 ();
 decap_12 FILLER_147_151 ();
 fill_4 FILLER_147_163 ();
 fill_1 FILLER_147_167 ();
 fill_4 FILLER_147_181 ();
 fill_1 FILLER_147_185 ();
 fill_2 FILLER_147_235 ();
 decap_12 FILLER_147_264 ();
 fill_4 FILLER_147_276 ();
 fill_2 FILLER_147_293 ();
 fill_2 FILLER_147_299 ();
 fill_1 FILLER_147_308 ();
 fill_1 FILLER_147_311 ();
 fill_2 FILLER_147_340 ();
 fill_2 FILLER_147_345 ();
 fill_1 FILLER_147_347 ();
 fill_1 FILLER_147_351 ();
 fill_2 FILLER_147_387 ();
 fill_1 FILLER_147_409 ();
 fill_2 FILLER_147_425 ();
 fill_1 FILLER_147_427 ();
 decap_12 FILLER_147_455 ();
 fill_2 FILLER_147_467 ();
 fill_2 FILLER_147_475 ();
 fill_2 FILLER_147_502 ();
 fill_4 FILLER_147_510 ();
 fill_1 FILLER_147_514 ();
 fill_2 FILLER_147_544 ();
 fill_1 FILLER_147_546 ();
 fill_4 FILLER_147_555 ();
 fill_1 FILLER_147_559 ();
 fill_8 FILLER_147_570 ();
 fill_2 FILLER_147_578 ();
 decap_12 FILLER_147_588 ();
 decap_12 FILLER_147_600 ();
 fill_4 FILLER_147_612 ();
 fill_2 FILLER_147_617 ();
 fill_4 FILLER_147_628 ();
 fill_1 FILLER_147_632 ();
 fill_2 FILLER_147_644 ();
 fill_1 FILLER_147_659 ();
 fill_1 FILLER_147_668 ();
 fill_2 FILLER_147_710 ();
 fill_4 FILLER_147_721 ();
 fill_2 FILLER_147_725 ();
 fill_1 FILLER_147_727 ();
 fill_1 FILLER_147_799 ();
 fill_1 FILLER_147_839 ();
 fill_1 FILLER_147_847 ();
 fill_1 FILLER_147_860 ();
 decap_12 FILLER_147_872 ();
 fill_1 FILLER_147_884 ();
 fill_8 FILLER_147_888 ();
 fill_4 FILLER_147_897 ();
 fill_1 FILLER_147_901 ();
 fill_4 FILLER_147_919 ();
 fill_1 FILLER_147_923 ();
 fill_4 FILLER_147_927 ();
 fill_2 FILLER_147_931 ();
 fill_1 FILLER_147_933 ();
 fill_2 FILLER_147_949 ();
 fill_1 FILLER_147_951 ();
 fill_4 FILLER_147_957 ();
 fill_2 FILLER_147_961 ();
 decap_12 FILLER_147_966 ();
 fill_2 FILLER_147_978 ();
 fill_1 FILLER_147_980 ();
 fill_4 FILLER_147_984 ();
 fill_4 FILLER_147_995 ();
 fill_2 FILLER_147_1012 ();
 fill_1 FILLER_147_1014 ();
 fill_8 FILLER_147_1027 ();
 fill_2 FILLER_147_1035 ();
 fill_1 FILLER_147_1037 ();
 decap_12 FILLER_148_3 ();
 decap_12 FILLER_148_15 ();
 fill_1 FILLER_148_27 ();
 fill_4 FILLER_148_29 ();
 fill_2 FILLER_148_33 ();
 fill_1 FILLER_148_35 ();
 fill_4 FILLER_148_56 ();
 fill_2 FILLER_148_60 ();
 fill_1 FILLER_148_62 ();
 fill_2 FILLER_148_81 ();
 fill_1 FILLER_148_83 ();
 fill_1 FILLER_148_85 ();
 fill_2 FILLER_148_104 ();
 fill_1 FILLER_148_106 ();
 fill_4 FILLER_148_136 ();
 fill_2 FILLER_148_141 ();
 fill_4 FILLER_148_152 ();
 fill_2 FILLER_148_156 ();
 fill_2 FILLER_148_178 ();
 fill_2 FILLER_148_194 ();
 fill_4 FILLER_148_235 ();
 fill_1 FILLER_148_239 ();
 fill_2 FILLER_148_263 ();
 fill_4 FILLER_148_336 ();
 fill_2 FILLER_148_340 ();
 fill_1 FILLER_148_342 ();
 fill_4 FILLER_148_414 ();
 fill_2 FILLER_148_418 ();
 fill_1 FILLER_148_421 ();
 fill_2 FILLER_148_427 ();
 fill_2 FILLER_148_439 ();
 decap_12 FILLER_148_444 ();
 fill_2 FILLER_148_456 ();
 fill_8 FILLER_148_461 ();
 fill_2 FILLER_148_469 ();
 fill_1 FILLER_148_475 ();
 fill_4 FILLER_148_477 ();
 fill_1 FILLER_148_481 ();
 fill_4 FILLER_148_502 ();
 fill_2 FILLER_148_529 ();
 fill_1 FILLER_148_531 ();
 fill_4 FILLER_148_555 ();
 fill_1 FILLER_148_559 ();
 fill_2 FILLER_148_576 ();
 fill_4 FILLER_148_583 ();
 fill_1 FILLER_148_587 ();
 fill_2 FILLER_148_589 ();
 fill_1 FILLER_148_606 ();
 fill_4 FILLER_148_613 ();
 fill_2 FILLER_148_617 ();
 fill_1 FILLER_148_619 ();
 fill_4 FILLER_148_628 ();
 fill_2 FILLER_148_632 ();
 fill_1 FILLER_148_634 ();
 fill_1 FILLER_148_643 ();
 fill_1 FILLER_148_648 ();
 fill_4 FILLER_148_670 ();
 fill_1 FILLER_148_674 ();
 fill_2 FILLER_148_698 ();
 fill_2 FILLER_148_715 ();
 fill_1 FILLER_148_717 ();
 fill_2 FILLER_148_805 ();
 fill_2 FILLER_148_847 ();
 fill_1 FILLER_148_849 ();
 fill_1 FILLER_148_863 ();
 fill_2 FILLER_148_869 ();
 fill_8 FILLER_148_884 ();
 fill_1 FILLER_148_892 ();
 fill_1 FILLER_148_904 ();
 fill_1 FILLER_148_931 ();
 fill_4 FILLER_148_973 ();
 fill_1 FILLER_148_1011 ();
 decap_12 FILLER_148_1019 ();
 fill_4 FILLER_148_1031 ();
 fill_1 FILLER_148_1035 ();
 fill_1 FILLER_148_1037 ();
 decap_12 FILLER_149_3 ();
 decap_12 FILLER_149_15 ();
 fill_4 FILLER_149_27 ();
 fill_2 FILLER_149_31 ();
 fill_1 FILLER_149_33 ();
 fill_2 FILLER_149_54 ();
 fill_2 FILLER_149_113 ();
 fill_2 FILLER_149_135 ();
 fill_8 FILLER_149_157 ();
 fill_2 FILLER_149_165 ();
 fill_1 FILLER_149_167 ();
 fill_2 FILLER_149_202 ();
 fill_1 FILLER_149_233 ();
 fill_1 FILLER_149_335 ();
 fill_1 FILLER_149_344 ();
 fill_1 FILLER_149_353 ();
 fill_1 FILLER_149_366 ();
 fill_1 FILLER_149_402 ();
 fill_2 FILLER_149_423 ();
 fill_1 FILLER_149_425 ();
 fill_1 FILLER_149_429 ();
 fill_1 FILLER_149_439 ();
 fill_4 FILLER_149_444 ();
 decap_12 FILLER_149_454 ();
 fill_2 FILLER_149_466 ();
 fill_8 FILLER_149_475 ();
 fill_2 FILLER_149_493 ();
 fill_4 FILLER_149_500 ();
 fill_4 FILLER_149_505 ();
 fill_1 FILLER_149_509 ();
 fill_2 FILLER_149_517 ();
 fill_1 FILLER_149_519 ();
 fill_4 FILLER_149_529 ();
 fill_1 FILLER_149_533 ();
 decap_12 FILLER_149_541 ();
 fill_4 FILLER_149_553 ();
 fill_2 FILLER_149_557 ();
 fill_1 FILLER_149_559 ();
 fill_2 FILLER_149_561 ();
 fill_4 FILLER_149_566 ();
 fill_1 FILLER_149_570 ();
 fill_1 FILLER_149_579 ();
 fill_8 FILLER_149_587 ();
 fill_1 FILLER_149_595 ();
 fill_1 FILLER_149_615 ();
 fill_2 FILLER_149_622 ();
 fill_2 FILLER_149_634 ();
 fill_1 FILLER_149_636 ();
 fill_4 FILLER_149_650 ();
 fill_1 FILLER_149_654 ();
 fill_4 FILLER_149_694 ();
 fill_2 FILLER_149_698 ();
 fill_1 FILLER_149_700 ();
 fill_4 FILLER_149_721 ();
 fill_2 FILLER_149_725 ();
 fill_1 FILLER_149_727 ();
 fill_2 FILLER_149_782 ();
 fill_2 FILLER_149_785 ();
 fill_1 FILLER_149_807 ();
 fill_2 FILLER_149_817 ();
 fill_4 FILLER_149_829 ();
 fill_4 FILLER_149_836 ();
 fill_4 FILLER_149_841 ();
 fill_4 FILLER_149_855 ();
 fill_2 FILLER_149_859 ();
 fill_1 FILLER_149_861 ();
 fill_4 FILLER_149_869 ();
 fill_2 FILLER_149_873 ();
 fill_2 FILLER_149_886 ();
 fill_1 FILLER_149_895 ();
 fill_1 FILLER_149_920 ();
 fill_1 FILLER_149_951 ();
 fill_2 FILLER_149_958 ();
 fill_2 FILLER_149_973 ();
 fill_8 FILLER_149_989 ();
 fill_2 FILLER_149_997 ();
 fill_4 FILLER_149_1002 ();
 fill_2 FILLER_149_1006 ();
 fill_4 FILLER_149_1009 ();
 fill_2 FILLER_149_1013 ();
 fill_2 FILLER_149_1035 ();
 fill_1 FILLER_149_1037 ();
 decap_12 FILLER_150_3 ();
 decap_12 FILLER_150_15 ();
 fill_1 FILLER_150_27 ();
 decap_12 FILLER_150_29 ();
 fill_2 FILLER_150_41 ();
 fill_2 FILLER_150_81 ();
 fill_1 FILLER_150_83 ();
 fill_4 FILLER_150_118 ();
 fill_1 FILLER_150_122 ();
 fill_2 FILLER_150_138 ();
 fill_2 FILLER_150_141 ();
 fill_1 FILLER_150_143 ();
 fill_2 FILLER_150_153 ();
 fill_2 FILLER_150_197 ();
 decap_12 FILLER_150_215 ();
 fill_1 FILLER_150_238 ();
 fill_4 FILLER_150_242 ();
 fill_2 FILLER_150_246 ();
 fill_2 FILLER_150_253 ();
 fill_1 FILLER_150_266 ();
 fill_1 FILLER_150_344 ();
 fill_2 FILLER_150_362 ();
 fill_2 FILLER_150_373 ();
 fill_2 FILLER_150_378 ();
 fill_1 FILLER_150_419 ();
 fill_1 FILLER_150_421 ();
 fill_1 FILLER_150_426 ();
 fill_1 FILLER_150_475 ();
 fill_4 FILLER_150_477 ();
 fill_1 FILLER_150_481 ();
 fill_4 FILLER_150_494 ();
 fill_2 FILLER_150_498 ();
 fill_2 FILLER_150_509 ();
 fill_4 FILLER_150_519 ();
 fill_2 FILLER_150_530 ();
 fill_1 FILLER_150_537 ();
 fill_1 FILLER_150_543 ();
 fill_4 FILLER_150_549 ();
 fill_2 FILLER_150_553 ();
 decap_12 FILLER_150_571 ();
 fill_4 FILLER_150_583 ();
 fill_1 FILLER_150_587 ();
 fill_2 FILLER_150_609 ();
 fill_1 FILLER_150_611 ();
 fill_4 FILLER_150_615 ();
 fill_2 FILLER_150_619 ();
 fill_2 FILLER_150_626 ();
 fill_4 FILLER_150_639 ();
 fill_1 FILLER_150_643 ();
 fill_4 FILLER_150_648 ();
 fill_1 FILLER_150_652 ();
 fill_1 FILLER_150_658 ();
 fill_4 FILLER_150_733 ();
 fill_2 FILLER_150_737 ();
 fill_1 FILLER_150_789 ();
 fill_2 FILLER_150_810 ();
 fill_1 FILLER_150_822 ();
 fill_1 FILLER_150_829 ();
 fill_4 FILLER_150_845 ();
 fill_1 FILLER_150_849 ();
 fill_2 FILLER_150_865 ();
 fill_1 FILLER_150_867 ();
 fill_2 FILLER_150_876 ();
 fill_1 FILLER_150_894 ();
 fill_8 FILLER_150_902 ();
 fill_1 FILLER_150_910 ();
 fill_1 FILLER_150_918 ();
 fill_1 FILLER_150_953 ();
 fill_2 FILLER_150_961 ();
 fill_4 FILLER_150_974 ();
 fill_2 FILLER_150_978 ();
 fill_8 FILLER_150_985 ();
 fill_1 FILLER_150_993 ();
 fill_2 FILLER_150_1010 ();
 fill_4 FILLER_150_1032 ();
 fill_1 FILLER_150_1037 ();
 decap_12 FILLER_151_3 ();
 decap_12 FILLER_151_15 ();
 fill_8 FILLER_151_27 ();
 fill_1 FILLER_151_35 ();
 fill_4 FILLER_151_66 ();
 fill_4 FILLER_151_99 ();
 fill_2 FILLER_151_113 ();
 fill_1 FILLER_151_115 ();
 fill_2 FILLER_151_156 ();
 fill_1 FILLER_151_158 ();
 fill_2 FILLER_151_178 ();
 fill_2 FILLER_151_225 ();
 fill_1 FILLER_151_235 ();
 fill_2 FILLER_151_268 ();
 fill_2 FILLER_151_291 ();
 fill_1 FILLER_151_335 ();
 fill_2 FILLER_151_362 ();
 fill_1 FILLER_151_375 ();
 fill_2 FILLER_151_379 ();
 fill_1 FILLER_151_381 ();
 fill_1 FILLER_151_388 ();
 fill_2 FILLER_151_393 ();
 fill_4 FILLER_151_403 ();
 fill_1 FILLER_151_407 ();
 fill_2 FILLER_151_436 ();
 fill_4 FILLER_151_444 ();
 fill_2 FILLER_151_456 ();
 fill_1 FILLER_151_503 ();
 fill_8 FILLER_151_505 ();
 fill_2 FILLER_151_513 ();
 fill_1 FILLER_151_515 ();
 fill_2 FILLER_151_526 ();
 fill_1 FILLER_151_528 ();
 fill_2 FILLER_151_534 ();
 fill_4 FILLER_151_547 ();
 fill_2 FILLER_151_551 ();
 fill_1 FILLER_151_592 ();
 fill_1 FILLER_151_615 ();
 fill_1 FILLER_151_617 ();
 fill_4 FILLER_151_664 ();
 fill_1 FILLER_151_668 ();
 fill_1 FILLER_151_673 ();
 fill_8 FILLER_151_720 ();
 fill_4 FILLER_151_802 ();
 fill_1 FILLER_151_806 ();
 fill_8 FILLER_151_823 ();
 fill_2 FILLER_151_831 ();
 fill_1 FILLER_151_833 ();
 fill_4 FILLER_151_845 ();
 fill_2 FILLER_151_950 ();
 fill_2 FILLER_151_1005 ();
 fill_1 FILLER_151_1007 ();
 decap_12 FILLER_151_1016 ();
 fill_8 FILLER_151_1028 ();
 fill_2 FILLER_151_1036 ();
 decap_12 FILLER_152_3 ();
 decap_12 FILLER_152_15 ();
 fill_1 FILLER_152_27 ();
 fill_4 FILLER_152_58 ();
 fill_1 FILLER_152_62 ();
 fill_1 FILLER_152_83 ();
 fill_4 FILLER_152_85 ();
 fill_1 FILLER_152_89 ();
 fill_1 FILLER_152_119 ();
 fill_2 FILLER_152_141 ();
 fill_4 FILLER_152_152 ();
 fill_2 FILLER_152_176 ();
 fill_2 FILLER_152_186 ();
 fill_1 FILLER_152_197 ();
 fill_1 FILLER_152_235 ();
 fill_1 FILLER_152_245 ();
 decap_12 FILLER_152_265 ();
 fill_1 FILLER_152_277 ();
 fill_1 FILLER_152_307 ();
 fill_2 FILLER_152_318 ();
 fill_1 FILLER_152_320 ();
 fill_2 FILLER_152_346 ();
 fill_4 FILLER_152_365 ();
 fill_2 FILLER_152_369 ();
 fill_1 FILLER_152_371 ();
 decap_12 FILLER_152_383 ();
 fill_4 FILLER_152_395 ();
 fill_2 FILLER_152_399 ();
 fill_1 FILLER_152_407 ();
 fill_2 FILLER_152_413 ();
 fill_1 FILLER_152_415 ();
 fill_1 FILLER_152_419 ();
 fill_4 FILLER_152_477 ();
 fill_2 FILLER_152_481 ();
 fill_1 FILLER_152_505 ();
 fill_1 FILLER_152_513 ();
 decap_12 FILLER_152_517 ();
 fill_2 FILLER_152_529 ();
 fill_1 FILLER_152_531 ();
 fill_2 FILLER_152_552 ();
 fill_1 FILLER_152_554 ();
 fill_1 FILLER_152_564 ();
 fill_4 FILLER_152_568 ();
 fill_8 FILLER_152_580 ();
 fill_4 FILLER_152_589 ();
 fill_8 FILLER_152_598 ();
 fill_2 FILLER_152_614 ();
 fill_1 FILLER_152_616 ();
 fill_1 FILLER_152_621 ();
 fill_4 FILLER_152_637 ();
 fill_2 FILLER_152_641 ();
 fill_1 FILLER_152_643 ();
 decap_12 FILLER_152_645 ();
 decap_12 FILLER_152_657 ();
 fill_4 FILLER_152_669 ();
 fill_2 FILLER_152_673 ();
 fill_8 FILLER_152_683 ();
 fill_4 FILLER_152_710 ();
 fill_1 FILLER_152_755 ();
 fill_1 FILLER_152_813 ();
 decap_12 FILLER_152_841 ();
 fill_2 FILLER_152_861 ();
 fill_2 FILLER_152_889 ();
 fill_1 FILLER_152_891 ();
 fill_8 FILLER_152_901 ();
 fill_1 FILLER_152_909 ();
 fill_2 FILLER_152_922 ();
 fill_2 FILLER_152_925 ();
 fill_4 FILLER_152_942 ();
 fill_2 FILLER_152_946 ();
 fill_1 FILLER_152_948 ();
 fill_4 FILLER_152_973 ();
 fill_2 FILLER_152_977 ();
 fill_1 FILLER_152_979 ();
 decap_12 FILLER_152_981 ();
 decap_12 FILLER_152_993 ();
 decap_12 FILLER_152_1005 ();
 decap_12 FILLER_152_1017 ();
 fill_4 FILLER_152_1029 ();
 fill_1 FILLER_152_1033 ();
 fill_1 FILLER_152_1037 ();
 decap_12 FILLER_153_3 ();
 decap_12 FILLER_153_15 ();
 fill_8 FILLER_153_27 ();
 fill_1 FILLER_153_35 ();
 fill_2 FILLER_153_57 ();
 fill_4 FILLER_153_108 ();
 fill_4 FILLER_153_113 ();
 fill_2 FILLER_153_117 ();
 fill_1 FILLER_153_119 ();
 fill_2 FILLER_153_140 ();
 fill_4 FILLER_153_162 ();
 fill_2 FILLER_153_166 ();
 fill_1 FILLER_153_169 ();
 fill_1 FILLER_153_190 ();
 fill_2 FILLER_153_215 ();
 fill_1 FILLER_153_217 ();
 fill_2 FILLER_153_225 ();
 fill_2 FILLER_153_241 ();
 fill_2 FILLER_153_251 ();
 fill_4 FILLER_153_267 ();
 fill_1 FILLER_153_279 ();
 fill_8 FILLER_153_281 ();
 fill_1 FILLER_153_289 ();
 fill_4 FILLER_153_299 ();
 fill_1 FILLER_153_327 ();
 fill_1 FILLER_153_337 ();
 fill_2 FILLER_153_374 ();
 fill_1 FILLER_153_384 ();
 decap_12 FILLER_153_413 ();
 fill_1 FILLER_153_425 ();
 fill_1 FILLER_153_435 ();
 fill_4 FILLER_153_443 ();
 fill_1 FILLER_153_447 ();
 fill_2 FILLER_153_475 ();
 fill_1 FILLER_153_491 ();
 fill_2 FILLER_153_501 ();
 fill_1 FILLER_153_503 ();
 decap_12 FILLER_153_505 ();
 decap_12 FILLER_153_517 ();
 decap_12 FILLER_153_529 ();
 fill_8 FILLER_153_541 ();
 fill_1 FILLER_153_549 ();
 fill_4 FILLER_153_555 ();
 fill_1 FILLER_153_559 ();
 fill_8 FILLER_153_567 ();
 fill_2 FILLER_153_575 ();
 fill_1 FILLER_153_577 ();
 fill_4 FILLER_153_586 ();
 fill_2 FILLER_153_590 ();
 fill_1 FILLER_153_592 ();
 decap_12 FILLER_153_600 ();
 fill_4 FILLER_153_612 ();
 fill_4 FILLER_153_622 ();
 fill_1 FILLER_153_626 ();
 decap_12 FILLER_153_634 ();
 decap_12 FILLER_153_646 ();
 fill_2 FILLER_153_658 ();
 fill_1 FILLER_153_660 ();
 fill_4 FILLER_153_666 ();
 fill_2 FILLER_153_670 ();
 fill_2 FILLER_153_681 ();
 fill_2 FILLER_153_726 ();
 fill_2 FILLER_153_729 ();
 fill_1 FILLER_153_731 ();
 fill_2 FILLER_153_761 ();
 fill_1 FILLER_153_763 ();
 fill_4 FILLER_153_780 ();
 fill_1 FILLER_153_785 ();
 decap_12 FILLER_153_795 ();
 fill_4 FILLER_153_807 ();
 fill_1 FILLER_153_811 ();
 fill_1 FILLER_153_872 ();
 fill_1 FILLER_153_889 ();
 fill_1 FILLER_153_895 ();
 fill_8 FILLER_153_900 ();
 fill_2 FILLER_153_908 ();
 fill_2 FILLER_153_915 ();
 fill_8 FILLER_153_922 ();
 fill_2 FILLER_153_939 ();
 fill_1 FILLER_153_944 ();
 fill_2 FILLER_153_950 ();
 fill_1 FILLER_153_957 ();
 decap_12 FILLER_153_980 ();
 decap_12 FILLER_153_992 ();
 fill_4 FILLER_153_1004 ();
 decap_12 FILLER_153_1009 ();
 fill_8 FILLER_153_1021 ();
 fill_2 FILLER_153_1029 ();
 fill_1 FILLER_153_1031 ();
 decap_12 FILLER_154_3 ();
 decap_12 FILLER_154_15 ();
 fill_1 FILLER_154_27 ();
 decap_12 FILLER_154_29 ();
 fill_2 FILLER_154_50 ();
 fill_2 FILLER_154_72 ();
 fill_1 FILLER_154_74 ();
 fill_4 FILLER_154_85 ();
 fill_2 FILLER_154_89 ();
 fill_1 FILLER_154_91 ();
 fill_1 FILLER_154_105 ();
 fill_4 FILLER_154_135 ();
 fill_1 FILLER_154_139 ();
 fill_4 FILLER_154_141 ();
 fill_1 FILLER_154_145 ();
 fill_4 FILLER_154_184 ();
 fill_2 FILLER_154_221 ();
 fill_1 FILLER_154_244 ();
 fill_1 FILLER_154_251 ();
 fill_1 FILLER_154_277 ();
 fill_1 FILLER_154_307 ();
 fill_1 FILLER_154_333 ();
 fill_4 FILLER_154_350 ();
 fill_2 FILLER_154_354 ();
 fill_2 FILLER_154_365 ();
 fill_1 FILLER_154_367 ();
 fill_4 FILLER_154_376 ();
 fill_2 FILLER_154_380 ();
 fill_2 FILLER_154_395 ();
 fill_2 FILLER_154_417 ();
 fill_1 FILLER_154_419 ();
 fill_2 FILLER_154_421 ();
 fill_8 FILLER_154_429 ();
 fill_2 FILLER_154_437 ();
 fill_8 FILLER_154_450 ();
 fill_2 FILLER_154_458 ();
 fill_1 FILLER_154_460 ();
 fill_4 FILLER_154_471 ();
 fill_1 FILLER_154_475 ();
 fill_4 FILLER_154_477 ();
 fill_1 FILLER_154_481 ();
 fill_1 FILLER_154_485 ();
 fill_4 FILLER_154_501 ();
 fill_1 FILLER_154_505 ();
 fill_4 FILLER_154_511 ();
 fill_2 FILLER_154_515 ();
 fill_1 FILLER_154_517 ();
 fill_4 FILLER_154_525 ();
 fill_2 FILLER_154_529 ();
 fill_1 FILLER_154_531 ();
 fill_8 FILLER_154_533 ();
 fill_2 FILLER_154_541 ();
 fill_2 FILLER_154_549 ();
 fill_1 FILLER_154_551 ();
 fill_8 FILLER_154_563 ();
 fill_8 FILLER_154_577 ();
 fill_2 FILLER_154_585 ();
 fill_1 FILLER_154_587 ();
 decap_12 FILLER_154_589 ();
 fill_4 FILLER_154_601 ();
 fill_8 FILLER_154_610 ();
 fill_8 FILLER_154_626 ();
 fill_2 FILLER_154_634 ();
 fill_1 FILLER_154_636 ();
 fill_1 FILLER_154_643 ();
 fill_4 FILLER_154_645 ();
 fill_2 FILLER_154_649 ();
 decap_12 FILLER_154_657 ();
 fill_4 FILLER_154_669 ();
 fill_2 FILLER_154_673 ();
 fill_4 FILLER_154_694 ();
 fill_2 FILLER_154_698 ();
 fill_2 FILLER_154_701 ();
 fill_1 FILLER_154_703 ();
 fill_2 FILLER_154_725 ();
 fill_1 FILLER_154_727 ();
 fill_2 FILLER_154_754 ();
 fill_1 FILLER_154_792 ();
 fill_1 FILLER_154_811 ();
 fill_1 FILLER_154_826 ();
 fill_2 FILLER_154_836 ();
 fill_4 FILLER_154_869 ();
 fill_1 FILLER_154_893 ();
 fill_1 FILLER_154_954 ();
 fill_4 FILLER_154_973 ();
 fill_2 FILLER_154_977 ();
 fill_1 FILLER_154_979 ();
 decap_12 FILLER_154_981 ();
 decap_12 FILLER_154_993 ();
 decap_12 FILLER_154_1005 ();
 decap_12 FILLER_154_1017 ();
 fill_4 FILLER_154_1029 ();
 fill_2 FILLER_154_1033 ();
 fill_1 FILLER_154_1035 ();
 fill_1 FILLER_154_1037 ();
 decap_12 FILLER_155_3 ();
 decap_12 FILLER_155_15 ();
 decap_12 FILLER_155_27 ();
 fill_2 FILLER_155_39 ();
 fill_1 FILLER_155_41 ();
 fill_4 FILLER_155_51 ();
 fill_1 FILLER_155_55 ();
 decap_12 FILLER_155_57 ();
 decap_12 FILLER_155_69 ();
 decap_12 FILLER_155_81 ();
 decap_12 FILLER_155_93 ();
 fill_4 FILLER_155_105 ();
 fill_2 FILLER_155_109 ();
 fill_1 FILLER_155_111 ();
 fill_1 FILLER_155_122 ();
 decap_12 FILLER_155_132 ();
 decap_12 FILLER_155_144 ();
 decap_12 FILLER_155_156 ();
 fill_2 FILLER_155_169 ();
 fill_2 FILLER_155_191 ();
 fill_2 FILLER_155_222 ();
 fill_2 FILLER_155_242 ();
 fill_2 FILLER_155_258 ();
 fill_4 FILLER_155_315 ();
 fill_1 FILLER_155_319 ();
 fill_4 FILLER_155_337 ();
 fill_2 FILLER_155_350 ();
 fill_4 FILLER_155_368 ();
 fill_4 FILLER_155_393 ();
 fill_2 FILLER_155_410 ();
 fill_2 FILLER_155_432 ();
 fill_8 FILLER_155_440 ();
 fill_4 FILLER_155_457 ();
 fill_2 FILLER_155_461 ();
 fill_1 FILLER_155_463 ();
 fill_2 FILLER_155_502 ();
 fill_8 FILLER_155_508 ();
 fill_1 FILLER_155_516 ();
 fill_8 FILLER_155_522 ();
 fill_2 FILLER_155_530 ();
 fill_8 FILLER_155_539 ();
 fill_2 FILLER_155_547 ();
 fill_1 FILLER_155_559 ();
 decap_12 FILLER_155_561 ();
 decap_12 FILLER_155_573 ();
 fill_4 FILLER_155_585 ();
 decap_12 FILLER_155_597 ();
 fill_4 FILLER_155_609 ();
 fill_2 FILLER_155_613 ();
 fill_1 FILLER_155_615 ();
 decap_12 FILLER_155_617 ();
 decap_12 FILLER_155_629 ();
 decap_12 FILLER_155_641 ();
 decap_12 FILLER_155_653 ();
 fill_4 FILLER_155_665 ();
 fill_2 FILLER_155_669 ();
 fill_1 FILLER_155_671 ();
 fill_8 FILLER_155_673 ();
 fill_1 FILLER_155_727 ();
 fill_2 FILLER_155_764 ();
 fill_1 FILLER_155_841 ();
 fill_4 FILLER_155_868 ();
 fill_1 FILLER_155_872 ();
 decap_12 FILLER_155_882 ();
 fill_2 FILLER_155_894 ();
 fill_1 FILLER_155_897 ();
 fill_2 FILLER_155_901 ();
 fill_4 FILLER_155_910 ();
 fill_2 FILLER_155_914 ();
 fill_8 FILLER_155_921 ();
 fill_1 FILLER_155_932 ();
 fill_2 FILLER_155_943 ();
 fill_4 FILLER_155_948 ();
 decap_12 FILLER_155_953 ();
 decap_12 FILLER_155_965 ();
 decap_12 FILLER_155_977 ();
 decap_12 FILLER_155_989 ();
 fill_4 FILLER_155_1001 ();
 fill_2 FILLER_155_1005 ();
 fill_1 FILLER_155_1007 ();
 decap_12 FILLER_155_1009 ();
 decap_12 FILLER_155_1021 ();
 fill_4 FILLER_155_1033 ();
 fill_1 FILLER_155_1037 ();
 decap_12 FILLER_156_3 ();
 decap_12 FILLER_156_15 ();
 fill_1 FILLER_156_27 ();
 decap_12 FILLER_156_29 ();
 decap_12 FILLER_156_41 ();
 decap_12 FILLER_156_53 ();
 decap_12 FILLER_156_65 ();
 fill_4 FILLER_156_77 ();
 fill_2 FILLER_156_81 ();
 fill_1 FILLER_156_83 ();
 decap_12 FILLER_156_85 ();
 decap_12 FILLER_156_97 ();
 decap_12 FILLER_156_109 ();
 decap_12 FILLER_156_121 ();
 fill_4 FILLER_156_133 ();
 fill_2 FILLER_156_137 ();
 fill_1 FILLER_156_139 ();
 decap_12 FILLER_156_141 ();
 decap_12 FILLER_156_153 ();
 fill_4 FILLER_156_165 ();
 fill_2 FILLER_156_169 ();
 fill_1 FILLER_156_171 ();
 fill_4 FILLER_156_192 ();
 fill_2 FILLER_156_197 ();
 fill_4 FILLER_156_210 ();
 fill_2 FILLER_156_250 ();
 fill_1 FILLER_156_263 ();
 fill_2 FILLER_156_267 ();
 fill_4 FILLER_156_276 ();
 fill_2 FILLER_156_280 ();
 fill_2 FILLER_156_306 ();
 fill_4 FILLER_156_318 ();
 fill_2 FILLER_156_421 ();
 fill_2 FILLER_156_427 ();
 fill_1 FILLER_156_441 ();
 decap_12 FILLER_156_448 ();
 fill_2 FILLER_156_467 ();
 fill_4 FILLER_156_472 ();
 fill_8 FILLER_156_477 ();
 fill_1 FILLER_156_485 ();
 fill_4 FILLER_156_499 ();
 fill_1 FILLER_156_503 ();
 fill_8 FILLER_156_524 ();
 decap_12 FILLER_156_533 ();
 fill_4 FILLER_156_560 ();
 fill_2 FILLER_156_573 ();
 fill_4 FILLER_156_582 ();
 fill_2 FILLER_156_586 ();
 fill_2 FILLER_156_589 ();
 fill_8 FILLER_156_596 ();
 fill_1 FILLER_156_604 ();
 decap_12 FILLER_156_610 ();
 decap_12 FILLER_156_622 ();
 fill_8 FILLER_156_634 ();
 fill_2 FILLER_156_642 ();
 decap_12 FILLER_156_645 ();
 decap_12 FILLER_156_657 ();
 fill_4 FILLER_156_669 ();
 fill_8 FILLER_156_678 ();
 fill_4 FILLER_156_701 ();
 fill_2 FILLER_156_729 ();
 fill_2 FILLER_156_753 ();
 fill_1 FILLER_156_755 ();
 fill_4 FILLER_156_805 ();
 fill_1 FILLER_156_869 ();
 decap_12 FILLER_156_890 ();
 decap_12 FILLER_156_902 ();
 fill_8 FILLER_156_914 ();
 fill_2 FILLER_156_922 ();
 decap_12 FILLER_156_925 ();
 decap_12 FILLER_156_937 ();
 decap_12 FILLER_156_949 ();
 decap_12 FILLER_156_961 ();
 fill_4 FILLER_156_973 ();
 fill_2 FILLER_156_977 ();
 fill_1 FILLER_156_979 ();
 decap_12 FILLER_156_981 ();
 decap_12 FILLER_156_993 ();
 decap_12 FILLER_156_1005 ();
 decap_12 FILLER_156_1017 ();
 fill_4 FILLER_156_1029 ();
 fill_2 FILLER_156_1033 ();
 fill_1 FILLER_156_1035 ();
 fill_1 FILLER_156_1037 ();
 decap_12 FILLER_157_5 ();
 decap_12 FILLER_157_17 ();
 decap_12 FILLER_157_29 ();
 decap_12 FILLER_157_41 ();
 fill_2 FILLER_157_53 ();
 fill_1 FILLER_157_55 ();
 decap_12 FILLER_157_57 ();
 decap_12 FILLER_157_69 ();
 decap_12 FILLER_157_81 ();
 decap_12 FILLER_157_93 ();
 fill_4 FILLER_157_105 ();
 fill_2 FILLER_157_109 ();
 fill_1 FILLER_157_111 ();
 decap_12 FILLER_157_113 ();
 decap_12 FILLER_157_125 ();
 decap_12 FILLER_157_137 ();
 decap_12 FILLER_157_149 ();
 fill_4 FILLER_157_161 ();
 fill_2 FILLER_157_165 ();
 fill_1 FILLER_157_167 ();
 fill_8 FILLER_157_169 ();
 fill_1 FILLER_157_177 ();
 fill_2 FILLER_157_189 ();
 fill_2 FILLER_157_219 ();
 fill_2 FILLER_157_225 ();
 fill_8 FILLER_157_245 ();
 fill_2 FILLER_157_253 ();
 fill_4 FILLER_157_281 ();
 fill_1 FILLER_157_285 ();
 fill_2 FILLER_157_295 ();
 fill_1 FILLER_157_317 ();
 fill_2 FILLER_157_326 ();
 fill_2 FILLER_157_341 ();
 fill_4 FILLER_157_355 ();
 fill_1 FILLER_157_359 ();
 fill_2 FILLER_157_407 ();
 fill_1 FILLER_157_409 ();
 fill_4 FILLER_157_442 ();
 fill_2 FILLER_157_446 ();
 decap_12 FILLER_157_449 ();
 fill_8 FILLER_157_461 ();
 fill_2 FILLER_157_469 ();
 fill_1 FILLER_157_483 ();
 fill_4 FILLER_157_489 ();
 fill_2 FILLER_157_501 ();
 fill_1 FILLER_157_503 ();
 decap_12 FILLER_157_505 ();
 fill_2 FILLER_157_517 ();
 fill_4 FILLER_157_525 ();
 fill_2 FILLER_157_529 ();
 fill_1 FILLER_157_531 ();
 fill_4 FILLER_157_539 ();
 fill_2 FILLER_157_558 ();
 decap_12 FILLER_157_568 ();
 decap_12 FILLER_157_580 ();
 fill_1 FILLER_157_592 ();
 decap_12 FILLER_157_598 ();
 fill_1 FILLER_157_610 ();
 fill_4 FILLER_157_617 ();
 fill_8 FILLER_157_628 ();
 fill_1 FILLER_157_636 ();
 decap_12 FILLER_157_643 ();
 fill_2 FILLER_157_655 ();
 fill_8 FILLER_157_663 ();
 fill_1 FILLER_157_671 ();
 fill_8 FILLER_157_673 ();
 fill_2 FILLER_157_701 ();
 fill_1 FILLER_157_703 ();
 fill_1 FILLER_157_742 ();
 fill_4 FILLER_157_785 ();
 fill_2 FILLER_157_789 ();
 decap_12 FILLER_157_802 ();
 decap_12 FILLER_157_814 ();
 fill_1 FILLER_157_826 ();
 fill_2 FILLER_157_830 ();
 fill_1 FILLER_157_832 ();
 fill_4 FILLER_157_836 ();
 fill_4 FILLER_157_869 ();
 fill_1 FILLER_157_873 ();
 decap_12 FILLER_157_879 ();
 fill_4 FILLER_157_891 ();
 fill_1 FILLER_157_895 ();
 decap_12 FILLER_157_897 ();
 decap_12 FILLER_157_909 ();
 decap_12 FILLER_157_921 ();
 decap_12 FILLER_157_933 ();
 fill_4 FILLER_157_945 ();
 fill_2 FILLER_157_949 ();
 fill_1 FILLER_157_951 ();
 decap_12 FILLER_157_953 ();
 decap_12 FILLER_157_965 ();
 decap_12 FILLER_157_977 ();
 decap_12 FILLER_157_989 ();
 fill_4 FILLER_157_1001 ();
 fill_2 FILLER_157_1005 ();
 fill_1 FILLER_157_1007 ();
 decap_12 FILLER_157_1009 ();
 decap_12 FILLER_157_1021 ();
 fill_4 FILLER_157_1033 ();
 fill_1 FILLER_157_1037 ();
 decap_12 FILLER_158_5 ();
 fill_8 FILLER_158_17 ();
 fill_2 FILLER_158_25 ();
 fill_1 FILLER_158_27 ();
 decap_12 FILLER_158_29 ();
 decap_12 FILLER_158_41 ();
 decap_12 FILLER_158_53 ();
 decap_12 FILLER_158_65 ();
 fill_4 FILLER_158_77 ();
 fill_2 FILLER_158_81 ();
 fill_1 FILLER_158_83 ();
 decap_12 FILLER_158_85 ();
 decap_12 FILLER_158_97 ();
 decap_12 FILLER_158_109 ();
 decap_12 FILLER_158_121 ();
 fill_4 FILLER_158_133 ();
 fill_2 FILLER_158_137 ();
 fill_1 FILLER_158_139 ();
 decap_12 FILLER_158_141 ();
 decap_12 FILLER_158_153 ();
 fill_4 FILLER_158_165 ();
 fill_1 FILLER_158_231 ();
 fill_4 FILLER_158_280 ();
 fill_2 FILLER_158_284 ();
 fill_1 FILLER_158_286 ();
 decap_12 FILLER_158_292 ();
 fill_4 FILLER_158_304 ();
 fill_2 FILLER_158_309 ();
 fill_1 FILLER_158_311 ();
 fill_1 FILLER_158_332 ();
 fill_1 FILLER_158_360 ();
 fill_1 FILLER_158_399 ();
 fill_4 FILLER_158_409 ();
 fill_2 FILLER_158_413 ();
 fill_1 FILLER_158_415 ();
 fill_2 FILLER_158_447 ();
 fill_1 FILLER_158_449 ();
 fill_4 FILLER_158_494 ();
 fill_2 FILLER_158_530 ();
 decap_12 FILLER_158_533 ();
 decap_12 FILLER_158_545 ();
 fill_4 FILLER_158_557 ();
 fill_2 FILLER_158_561 ();
 fill_1 FILLER_158_563 ();
 fill_2 FILLER_158_570 ();
 fill_1 FILLER_158_572 ();
 fill_1 FILLER_158_576 ();
 fill_1 FILLER_158_587 ();
 fill_2 FILLER_158_589 ();
 decap_12 FILLER_158_618 ();
 decap_12 FILLER_158_630 ();
 fill_2 FILLER_158_642 ();
 decap_12 FILLER_158_645 ();
 decap_12 FILLER_158_657 ();
 decap_12 FILLER_158_669 ();
 fill_1 FILLER_158_699 ();
 fill_2 FILLER_158_744 ();
 fill_1 FILLER_158_746 ();
 fill_4 FILLER_158_752 ();
 fill_4 FILLER_158_803 ();
 fill_1 FILLER_158_807 ();
 fill_1 FILLER_158_811 ();
 fill_2 FILLER_158_821 ();
 fill_1 FILLER_158_823 ();
 fill_2 FILLER_158_836 ();
 fill_1 FILLER_158_867 ();
 fill_1 FILLER_158_869 ();
 decap_12 FILLER_158_886 ();
 decap_12 FILLER_158_898 ();
 decap_12 FILLER_158_910 ();
 fill_2 FILLER_158_922 ();
 decap_12 FILLER_158_925 ();
 decap_12 FILLER_158_937 ();
 decap_12 FILLER_158_949 ();
 decap_12 FILLER_158_961 ();
 fill_4 FILLER_158_973 ();
 fill_2 FILLER_158_977 ();
 fill_1 FILLER_158_979 ();
 decap_12 FILLER_158_981 ();
 decap_12 FILLER_158_993 ();
 decap_12 FILLER_158_1005 ();
 decap_12 FILLER_158_1017 ();
 fill_4 FILLER_158_1029 ();
 fill_2 FILLER_158_1033 ();
 fill_1 FILLER_158_1035 ();
 fill_1 FILLER_158_1037 ();
 decap_12 FILLER_159_5 ();
 decap_12 FILLER_159_17 ();
 decap_12 FILLER_159_29 ();
 decap_12 FILLER_159_41 ();
 fill_2 FILLER_159_53 ();
 fill_1 FILLER_159_55 ();
 decap_12 FILLER_159_57 ();
 decap_12 FILLER_159_69 ();
 decap_12 FILLER_159_81 ();
 decap_12 FILLER_159_93 ();
 fill_4 FILLER_159_105 ();
 fill_2 FILLER_159_109 ();
 fill_1 FILLER_159_111 ();
 decap_12 FILLER_159_113 ();
 decap_12 FILLER_159_125 ();
 decap_12 FILLER_159_137 ();
 decap_12 FILLER_159_149 ();
 fill_4 FILLER_159_161 ();
 fill_2 FILLER_159_165 ();
 fill_1 FILLER_159_167 ();
 fill_4 FILLER_159_206 ();
 fill_4 FILLER_159_218 ();
 fill_2 FILLER_159_222 ();
 fill_2 FILLER_159_254 ();
 fill_1 FILLER_159_256 ();
 fill_2 FILLER_159_297 ();
 fill_4 FILLER_159_308 ();
 fill_1 FILLER_159_312 ();
 fill_2 FILLER_159_345 ();
 fill_1 FILLER_159_347 ();
 fill_4 FILLER_159_362 ();
 fill_2 FILLER_159_366 ();
 fill_1 FILLER_159_368 ();
 fill_2 FILLER_159_389 ();
 fill_1 FILLER_159_391 ();
 fill_2 FILLER_159_402 ();
 fill_1 FILLER_159_404 ();
 fill_2 FILLER_159_446 ();
 fill_2 FILLER_159_449 ();
 fill_1 FILLER_159_459 ();
 fill_1 FILLER_159_476 ();
 fill_1 FILLER_159_490 ();
 fill_1 FILLER_159_503 ();
 fill_1 FILLER_159_505 ();
 fill_4 FILLER_159_511 ();
 fill_2 FILLER_159_515 ();
 fill_4 FILLER_159_520 ();
 fill_4 FILLER_159_531 ();
 fill_2 FILLER_159_585 ();
 fill_1 FILLER_159_587 ();
 fill_2 FILLER_159_600 ();
 fill_4 FILLER_159_610 ();
 fill_2 FILLER_159_614 ();
 fill_4 FILLER_159_622 ();
 fill_2 FILLER_159_626 ();
 decap_12 FILLER_159_643 ();
 fill_4 FILLER_159_655 ();
 fill_2 FILLER_159_659 ();
 fill_2 FILLER_159_669 ();
 fill_1 FILLER_159_671 ();
 fill_8 FILLER_159_673 ();
 fill_1 FILLER_159_681 ();
 fill_1 FILLER_159_690 ();
 decap_12 FILLER_159_707 ();
 fill_4 FILLER_159_722 ();
 fill_2 FILLER_159_726 ();
 fill_8 FILLER_159_729 ();
 fill_2 FILLER_159_737 ();
 fill_8 FILLER_159_760 ();
 fill_1 FILLER_159_768 ();
 fill_1 FILLER_159_821 ();
 fill_2 FILLER_159_838 ();
 fill_4 FILLER_159_850 ();
 fill_2 FILLER_159_854 ();
 fill_1 FILLER_159_856 ();
 fill_2 FILLER_159_866 ();
 fill_1 FILLER_159_868 ();
 fill_4 FILLER_159_891 ();
 fill_1 FILLER_159_895 ();
 decap_12 FILLER_159_897 ();
 decap_12 FILLER_159_909 ();
 decap_12 FILLER_159_921 ();
 decap_12 FILLER_159_933 ();
 fill_4 FILLER_159_945 ();
 fill_2 FILLER_159_949 ();
 fill_1 FILLER_159_951 ();
 decap_12 FILLER_159_953 ();
 decap_12 FILLER_159_965 ();
 decap_12 FILLER_159_977 ();
 decap_12 FILLER_159_989 ();
 fill_4 FILLER_159_1001 ();
 fill_2 FILLER_159_1005 ();
 fill_1 FILLER_159_1007 ();
 decap_12 FILLER_159_1009 ();
 decap_12 FILLER_159_1021 ();
 fill_4 FILLER_159_1033 ();
 fill_1 FILLER_159_1037 ();
 decap_12 FILLER_160_5 ();
 fill_8 FILLER_160_17 ();
 fill_2 FILLER_160_25 ();
 fill_1 FILLER_160_27 ();
 decap_12 FILLER_160_29 ();
 decap_12 FILLER_160_41 ();
 decap_12 FILLER_160_53 ();
 decap_12 FILLER_160_65 ();
 fill_4 FILLER_160_77 ();
 fill_2 FILLER_160_81 ();
 fill_1 FILLER_160_83 ();
 decap_12 FILLER_160_85 ();
 decap_12 FILLER_160_97 ();
 decap_12 FILLER_160_109 ();
 decap_12 FILLER_160_121 ();
 fill_4 FILLER_160_133 ();
 fill_2 FILLER_160_137 ();
 fill_1 FILLER_160_139 ();
 decap_12 FILLER_160_141 ();
 decap_12 FILLER_160_153 ();
 decap_12 FILLER_160_165 ();
 decap_12 FILLER_160_177 ();
 fill_1 FILLER_160_189 ();
 fill_2 FILLER_160_193 ();
 fill_1 FILLER_160_195 ();
 decap_12 FILLER_160_197 ();
 fill_2 FILLER_160_209 ();
 fill_1 FILLER_160_211 ();
 fill_1 FILLER_160_262 ();
 fill_1 FILLER_160_275 ();
 fill_1 FILLER_160_309 ();
 fill_4 FILLER_160_350 ();
 fill_1 FILLER_160_354 ();
 fill_4 FILLER_160_370 ();
 fill_2 FILLER_160_410 ();
 fill_2 FILLER_160_418 ();
 fill_2 FILLER_160_421 ();
 fill_2 FILLER_160_447 ();
 fill_1 FILLER_160_475 ();
 fill_4 FILLER_160_500 ();
 fill_2 FILLER_160_504 ();
 fill_1 FILLER_160_506 ();
 fill_1 FILLER_160_510 ();
 decap_12 FILLER_160_518 ();
 fill_2 FILLER_160_530 ();
 decap_12 FILLER_160_533 ();
 decap_12 FILLER_160_545 ();
 fill_4 FILLER_160_557 ();
 fill_1 FILLER_160_561 ();
 decap_12 FILLER_160_574 ();
 fill_2 FILLER_160_586 ();
 fill_4 FILLER_160_589 ();
 fill_2 FILLER_160_593 ();
 fill_1 FILLER_160_595 ();
 decap_12 FILLER_160_604 ();
 fill_8 FILLER_160_616 ();
 fill_2 FILLER_160_624 ();
 fill_4 FILLER_160_632 ();
 fill_1 FILLER_160_636 ();
 fill_2 FILLER_160_641 ();
 fill_1 FILLER_160_643 ();
 fill_2 FILLER_160_645 ();
 fill_1 FILLER_160_647 ();
 decap_12 FILLER_160_654 ();
 fill_8 FILLER_160_672 ();
 fill_2 FILLER_160_680 ();
 fill_2 FILLER_160_698 ();
 fill_1 FILLER_160_709 ();
 fill_2 FILLER_160_729 ();
 fill_1 FILLER_160_731 ();
 fill_4 FILLER_160_757 ();
 fill_2 FILLER_160_761 ();
 fill_2 FILLER_160_768 ();
 fill_2 FILLER_160_780 ();
 fill_4 FILLER_160_787 ();
 fill_2 FILLER_160_791 ();
 fill_2 FILLER_160_810 ();
 fill_1 FILLER_160_818 ();
 fill_2 FILLER_160_827 ();
 fill_2 FILLER_160_837 ();
 fill_1 FILLER_160_839 ();
 fill_2 FILLER_160_866 ();
 decap_12 FILLER_160_888 ();
 decap_12 FILLER_160_900 ();
 decap_12 FILLER_160_912 ();
 decap_12 FILLER_160_925 ();
 decap_12 FILLER_160_937 ();
 decap_12 FILLER_160_949 ();
 decap_12 FILLER_160_961 ();
 fill_4 FILLER_160_973 ();
 fill_2 FILLER_160_977 ();
 fill_1 FILLER_160_979 ();
 decap_12 FILLER_160_981 ();
 decap_12 FILLER_160_993 ();
 decap_12 FILLER_160_1005 ();
 decap_12 FILLER_160_1017 ();
 fill_4 FILLER_160_1029 ();
 fill_2 FILLER_160_1033 ();
 fill_1 FILLER_160_1035 ();
 fill_1 FILLER_160_1037 ();
 decap_12 FILLER_161_5 ();
 decap_12 FILLER_161_17 ();
 decap_12 FILLER_161_29 ();
 decap_12 FILLER_161_41 ();
 fill_2 FILLER_161_53 ();
 fill_1 FILLER_161_55 ();
 decap_12 FILLER_161_57 ();
 decap_12 FILLER_161_69 ();
 decap_12 FILLER_161_81 ();
 decap_12 FILLER_161_93 ();
 fill_4 FILLER_161_105 ();
 fill_2 FILLER_161_109 ();
 fill_1 FILLER_161_111 ();
 decap_12 FILLER_161_113 ();
 decap_12 FILLER_161_125 ();
 decap_12 FILLER_161_137 ();
 decap_12 FILLER_161_149 ();
 fill_4 FILLER_161_161 ();
 fill_2 FILLER_161_165 ();
 fill_1 FILLER_161_167 ();
 decap_12 FILLER_161_169 ();
 decap_12 FILLER_161_181 ();
 decap_12 FILLER_161_193 ();
 decap_12 FILLER_161_205 ();
 fill_4 FILLER_161_217 ();
 fill_2 FILLER_161_221 ();
 fill_1 FILLER_161_223 ();
 fill_1 FILLER_161_225 ();
 fill_4 FILLER_161_235 ();
 fill_2 FILLER_161_239 ();
 fill_8 FILLER_161_250 ();
 fill_2 FILLER_161_258 ();
 fill_4 FILLER_161_267 ();
 fill_1 FILLER_161_279 ();
 fill_1 FILLER_161_288 ();
 fill_2 FILLER_161_296 ();
 fill_2 FILLER_161_334 ();
 fill_4 FILLER_161_337 ();
 fill_2 FILLER_161_389 ();
 fill_1 FILLER_161_391 ();
 fill_1 FILLER_161_435 ();
 fill_2 FILLER_161_445 ();
 fill_1 FILLER_161_447 ();
 fill_2 FILLER_161_456 ();
 fill_1 FILLER_161_458 ();
 fill_2 FILLER_161_474 ();
 fill_1 FILLER_161_476 ();
 fill_2 FILLER_161_484 ();
 fill_1 FILLER_161_497 ();
 fill_1 FILLER_161_503 ();
 fill_8 FILLER_161_509 ();
 decap_12 FILLER_161_520 ();
 decap_12 FILLER_161_532 ();
 fill_8 FILLER_161_544 ();
 fill_2 FILLER_161_552 ();
 fill_1 FILLER_161_554 ();
 fill_4 FILLER_161_574 ();
 fill_1 FILLER_161_578 ();
 fill_8 FILLER_161_586 ();
 fill_2 FILLER_161_594 ();
 decap_12 FILLER_161_602 ();
 fill_2 FILLER_161_614 ();
 decap_12 FILLER_161_617 ();
 decap_12 FILLER_161_629 ();
 fill_4 FILLER_161_641 ();
 fill_1 FILLER_161_645 ();
 decap_12 FILLER_161_651 ();
 fill_8 FILLER_161_663 ();
 fill_1 FILLER_161_671 ();
 fill_8 FILLER_161_673 ();
 fill_4 FILLER_161_684 ();
 fill_2 FILLER_161_688 ();
 fill_4 FILLER_161_723 ();
 fill_1 FILLER_161_727 ();
 fill_1 FILLER_161_729 ();
 fill_2 FILLER_161_768 ();
 fill_1 FILLER_161_785 ();
 fill_4 FILLER_161_823 ();
 fill_2 FILLER_161_827 ();
 fill_1 FILLER_161_829 ();
 fill_2 FILLER_161_837 ();
 fill_1 FILLER_161_839 ();
 decap_12 FILLER_161_841 ();
 decap_12 FILLER_161_853 ();
 fill_4 FILLER_161_865 ();
 fill_2 FILLER_161_869 ();
 fill_1 FILLER_161_871 ();
 decap_12 FILLER_161_878 ();
 fill_4 FILLER_161_890 ();
 fill_2 FILLER_161_894 ();
 decap_12 FILLER_161_897 ();
 decap_12 FILLER_161_909 ();
 decap_12 FILLER_161_921 ();
 decap_12 FILLER_161_933 ();
 fill_4 FILLER_161_945 ();
 fill_2 FILLER_161_949 ();
 fill_1 FILLER_161_951 ();
 decap_12 FILLER_161_953 ();
 decap_12 FILLER_161_965 ();
 decap_12 FILLER_161_977 ();
 decap_12 FILLER_161_989 ();
 fill_4 FILLER_161_1001 ();
 fill_2 FILLER_161_1005 ();
 fill_1 FILLER_161_1007 ();
 decap_12 FILLER_161_1009 ();
 decap_12 FILLER_161_1021 ();
 fill_4 FILLER_161_1033 ();
 fill_1 FILLER_161_1037 ();
 decap_12 FILLER_162_7 ();
 fill_8 FILLER_162_19 ();
 fill_1 FILLER_162_27 ();
 decap_12 FILLER_162_29 ();
 decap_12 FILLER_162_41 ();
 decap_12 FILLER_162_53 ();
 decap_12 FILLER_162_65 ();
 fill_4 FILLER_162_77 ();
 fill_2 FILLER_162_81 ();
 fill_1 FILLER_162_83 ();
 decap_12 FILLER_162_85 ();
 decap_12 FILLER_162_97 ();
 decap_12 FILLER_162_109 ();
 decap_12 FILLER_162_121 ();
 fill_4 FILLER_162_133 ();
 fill_2 FILLER_162_137 ();
 fill_1 FILLER_162_139 ();
 decap_12 FILLER_162_141 ();
 decap_12 FILLER_162_153 ();
 decap_12 FILLER_162_165 ();
 decap_12 FILLER_162_177 ();
 fill_4 FILLER_162_189 ();
 fill_2 FILLER_162_193 ();
 fill_1 FILLER_162_195 ();
 decap_12 FILLER_162_197 ();
 decap_12 FILLER_162_209 ();
 fill_2 FILLER_162_221 ();
 fill_4 FILLER_162_253 ();
 fill_1 FILLER_162_257 ();
 fill_1 FILLER_162_300 ();
 fill_1 FILLER_162_312 ();
 fill_4 FILLER_162_334 ();
 decap_12 FILLER_162_343 ();
 fill_4 FILLER_162_359 ();
 fill_1 FILLER_162_363 ();
 fill_2 FILLER_162_365 ();
 fill_2 FILLER_162_372 ();
 decap_12 FILLER_162_382 ();
 fill_1 FILLER_162_394 ();
 fill_2 FILLER_162_428 ();
 fill_2 FILLER_162_474 ();
 fill_4 FILLER_162_477 ();
 fill_2 FILLER_162_494 ();
 fill_2 FILLER_162_504 ();
 fill_1 FILLER_162_506 ();
 fill_8 FILLER_162_515 ();
 fill_4 FILLER_162_526 ();
 fill_2 FILLER_162_530 ();
 decap_12 FILLER_162_548 ();
 fill_2 FILLER_162_560 ();
 fill_1 FILLER_162_562 ();
 decap_12 FILLER_162_575 ();
 fill_1 FILLER_162_587 ();
 decap_12 FILLER_162_589 ();
 fill_8 FILLER_162_601 ();
 decap_12 FILLER_162_614 ();
 decap_12 FILLER_162_626 ();
 fill_4 FILLER_162_638 ();
 fill_2 FILLER_162_642 ();
 decap_12 FILLER_162_645 ();
 fill_8 FILLER_162_657 ();
 fill_2 FILLER_162_665 ();
 fill_2 FILLER_162_698 ();
 fill_1 FILLER_162_709 ();
 fill_2 FILLER_162_713 ();
 fill_1 FILLER_162_755 ();
 fill_4 FILLER_162_757 ();
 fill_2 FILLER_162_761 ();
 fill_2 FILLER_162_778 ();
 fill_2 FILLER_162_786 ();
 fill_4 FILLER_162_805 ();
 fill_2 FILLER_162_809 ();
 fill_1 FILLER_162_811 ();
 fill_1 FILLER_162_830 ();
 fill_1 FILLER_162_867 ();
 decap_12 FILLER_162_895 ();
 decap_12 FILLER_162_907 ();
 fill_4 FILLER_162_919 ();
 fill_1 FILLER_162_923 ();
 decap_12 FILLER_162_925 ();
 decap_12 FILLER_162_937 ();
 decap_12 FILLER_162_949 ();
 decap_12 FILLER_162_961 ();
 fill_4 FILLER_162_973 ();
 fill_2 FILLER_162_977 ();
 fill_1 FILLER_162_979 ();
 decap_12 FILLER_162_981 ();
 decap_12 FILLER_162_993 ();
 decap_12 FILLER_162_1005 ();
 decap_12 FILLER_162_1017 ();
 fill_1 FILLER_162_1029 ();
 fill_1 FILLER_162_1037 ();
 decap_12 FILLER_163_5 ();
 decap_12 FILLER_163_17 ();
 decap_12 FILLER_163_29 ();
 decap_12 FILLER_163_41 ();
 fill_2 FILLER_163_53 ();
 fill_1 FILLER_163_55 ();
 decap_12 FILLER_163_57 ();
 decap_12 FILLER_163_69 ();
 decap_12 FILLER_163_81 ();
 decap_12 FILLER_163_93 ();
 fill_4 FILLER_163_105 ();
 fill_2 FILLER_163_109 ();
 fill_1 FILLER_163_111 ();
 decap_12 FILLER_163_113 ();
 decap_12 FILLER_163_125 ();
 decap_12 FILLER_163_137 ();
 decap_12 FILLER_163_149 ();
 fill_4 FILLER_163_161 ();
 fill_2 FILLER_163_165 ();
 fill_1 FILLER_163_167 ();
 decap_12 FILLER_163_169 ();
 decap_12 FILLER_163_181 ();
 decap_12 FILLER_163_193 ();
 decap_12 FILLER_163_205 ();
 fill_4 FILLER_163_217 ();
 fill_2 FILLER_163_221 ();
 fill_1 FILLER_163_223 ();
 decap_12 FILLER_163_245 ();
 fill_4 FILLER_163_257 ();
 fill_1 FILLER_163_261 ();
 fill_1 FILLER_163_266 ();
 fill_4 FILLER_163_275 ();
 fill_1 FILLER_163_279 ();
 fill_2 FILLER_163_289 ();
 fill_1 FILLER_163_302 ();
 fill_4 FILLER_163_307 ();
 fill_1 FILLER_163_332 ();
 fill_1 FILLER_163_358 ();
 fill_4 FILLER_163_386 ();
 fill_2 FILLER_163_390 ();
 fill_1 FILLER_163_416 ();
 fill_2 FILLER_163_446 ();
 fill_2 FILLER_163_458 ();
 fill_2 FILLER_163_474 ();
 fill_4 FILLER_163_482 ();
 fill_1 FILLER_163_489 ();
 fill_4 FILLER_163_499 ();
 fill_1 FILLER_163_503 ();
 fill_2 FILLER_163_505 ();
 decap_12 FILLER_163_515 ();
 decap_12 FILLER_163_527 ();
 decap_12 FILLER_163_539 ();
 fill_8 FILLER_163_551 ();
 fill_1 FILLER_163_559 ();
 decap_12 FILLER_163_561 ();
 decap_12 FILLER_163_573 ();
 fill_8 FILLER_163_585 ();
 fill_2 FILLER_163_593 ();
 decap_12 FILLER_163_601 ();
 fill_2 FILLER_163_613 ();
 fill_1 FILLER_163_615 ();
 fill_8 FILLER_163_617 ();
 fill_1 FILLER_163_625 ();
 decap_12 FILLER_163_632 ();
 decap_12 FILLER_163_644 ();
 fill_4 FILLER_163_656 ();
 fill_2 FILLER_163_660 ();
 fill_4 FILLER_163_667 ();
 fill_1 FILLER_163_671 ();
 decap_12 FILLER_163_673 ();
 decap_12 FILLER_163_685 ();
 decap_12 FILLER_163_697 ();
 decap_12 FILLER_163_709 ();
 fill_4 FILLER_163_721 ();
 fill_2 FILLER_163_725 ();
 fill_1 FILLER_163_727 ();
 fill_1 FILLER_163_738 ();
 fill_2 FILLER_163_758 ();
 fill_4 FILLER_163_779 ();
 fill_1 FILLER_163_783 ();
 fill_1 FILLER_163_799 ();
 fill_4 FILLER_163_808 ();
 fill_2 FILLER_163_812 ();
 fill_8 FILLER_163_822 ();
 fill_1 FILLER_163_830 ();
 fill_1 FILLER_163_839 ();
 fill_1 FILLER_163_841 ();
 fill_4 FILLER_163_869 ();
 fill_1 FILLER_163_873 ();
 fill_2 FILLER_163_880 ();
 fill_1 FILLER_163_882 ();
 fill_2 FILLER_163_894 ();
 decap_12 FILLER_163_902 ();
 decap_12 FILLER_163_914 ();
 decap_12 FILLER_163_926 ();
 decap_12 FILLER_163_938 ();
 fill_2 FILLER_163_950 ();
 decap_12 FILLER_163_953 ();
 decap_12 FILLER_163_965 ();
 decap_12 FILLER_163_977 ();
 decap_12 FILLER_163_989 ();
 fill_4 FILLER_163_1001 ();
 fill_2 FILLER_163_1005 ();
 fill_1 FILLER_163_1007 ();
 decap_12 FILLER_163_1009 ();
 decap_12 FILLER_163_1021 ();
 fill_4 FILLER_163_1033 ();
 fill_1 FILLER_163_1037 ();
 decap_12 FILLER_164_5 ();
 fill_8 FILLER_164_17 ();
 fill_2 FILLER_164_25 ();
 fill_1 FILLER_164_27 ();
 decap_12 FILLER_164_29 ();
 decap_12 FILLER_164_41 ();
 decap_12 FILLER_164_53 ();
 decap_12 FILLER_164_65 ();
 fill_4 FILLER_164_77 ();
 fill_2 FILLER_164_81 ();
 fill_1 FILLER_164_83 ();
 decap_12 FILLER_164_85 ();
 decap_12 FILLER_164_97 ();
 decap_12 FILLER_164_109 ();
 decap_12 FILLER_164_121 ();
 fill_4 FILLER_164_133 ();
 fill_2 FILLER_164_137 ();
 fill_1 FILLER_164_139 ();
 decap_12 FILLER_164_141 ();
 decap_12 FILLER_164_153 ();
 decap_12 FILLER_164_165 ();
 decap_12 FILLER_164_177 ();
 fill_4 FILLER_164_189 ();
 fill_2 FILLER_164_193 ();
 fill_1 FILLER_164_195 ();
 decap_12 FILLER_164_197 ();
 decap_12 FILLER_164_209 ();
 fill_8 FILLER_164_221 ();
 fill_2 FILLER_164_229 ();
 fill_8 FILLER_164_261 ();
 fill_4 FILLER_164_272 ();
 fill_2 FILLER_164_276 ();
 fill_1 FILLER_164_278 ();
 fill_1 FILLER_164_284 ();
 fill_4 FILLER_164_309 ();
 fill_2 FILLER_164_313 ();
 fill_2 FILLER_164_329 ();
 fill_1 FILLER_164_374 ();
 fill_1 FILLER_164_387 ();
 fill_2 FILLER_164_418 ();
 fill_8 FILLER_164_507 ();
 fill_1 FILLER_164_515 ();
 fill_8 FILLER_164_521 ();
 fill_2 FILLER_164_529 ();
 fill_1 FILLER_164_531 ();
 decap_12 FILLER_164_533 ();
 fill_2 FILLER_164_545 ();
 fill_1 FILLER_164_547 ();
 fill_4 FILLER_164_556 ();
 fill_1 FILLER_164_560 ();
 fill_2 FILLER_164_567 ();
 fill_4 FILLER_164_574 ();
 fill_2 FILLER_164_578 ();
 fill_1 FILLER_164_580 ();
 fill_2 FILLER_164_586 ();
 decap_12 FILLER_164_589 ();
 decap_12 FILLER_164_601 ();
 decap_12 FILLER_164_613 ();
 decap_12 FILLER_164_625 ();
 fill_4 FILLER_164_637 ();
 fill_2 FILLER_164_641 ();
 fill_1 FILLER_164_643 ();
 decap_12 FILLER_164_651 ();
 fill_8 FILLER_164_663 ();
 decap_12 FILLER_164_687 ();
 fill_1 FILLER_164_699 ();
 decap_12 FILLER_164_701 ();
 decap_12 FILLER_164_713 ();
 fill_4 FILLER_164_725 ();
 fill_2 FILLER_164_729 ();
 fill_2 FILLER_164_734 ();
 fill_1 FILLER_164_736 ();
 fill_4 FILLER_164_760 ();
 fill_8 FILLER_164_767 ();
 decap_12 FILLER_164_782 ();
 fill_1 FILLER_164_794 ();
 fill_1 FILLER_164_811 ();
 fill_1 FILLER_164_813 ();
 fill_2 FILLER_164_832 ();
 fill_8 FILLER_164_854 ();
 fill_2 FILLER_164_865 ();
 fill_1 FILLER_164_867 ();
 fill_1 FILLER_164_882 ();
 decap_12 FILLER_164_896 ();
 decap_12 FILLER_164_908 ();
 fill_4 FILLER_164_920 ();
 decap_12 FILLER_164_925 ();
 decap_12 FILLER_164_937 ();
 decap_12 FILLER_164_949 ();
 decap_12 FILLER_164_961 ();
 fill_4 FILLER_164_973 ();
 fill_2 FILLER_164_977 ();
 fill_1 FILLER_164_979 ();
 decap_12 FILLER_164_981 ();
 decap_12 FILLER_164_993 ();
 decap_12 FILLER_164_1005 ();
 decap_12 FILLER_164_1017 ();
 fill_4 FILLER_164_1029 ();
 fill_2 FILLER_164_1033 ();
 fill_1 FILLER_164_1035 ();
 fill_1 FILLER_164_1037 ();
 decap_12 FILLER_165_5 ();
 decap_12 FILLER_165_17 ();
 decap_12 FILLER_165_29 ();
 decap_12 FILLER_165_41 ();
 fill_2 FILLER_165_53 ();
 fill_1 FILLER_165_55 ();
 decap_12 FILLER_165_57 ();
 decap_12 FILLER_165_69 ();
 decap_12 FILLER_165_81 ();
 decap_12 FILLER_165_93 ();
 fill_4 FILLER_165_105 ();
 fill_2 FILLER_165_109 ();
 fill_1 FILLER_165_111 ();
 decap_12 FILLER_165_113 ();
 decap_12 FILLER_165_125 ();
 decap_12 FILLER_165_137 ();
 decap_12 FILLER_165_149 ();
 fill_4 FILLER_165_161 ();
 fill_2 FILLER_165_165 ();
 fill_1 FILLER_165_167 ();
 decap_12 FILLER_165_169 ();
 decap_12 FILLER_165_181 ();
 decap_12 FILLER_165_193 ();
 decap_12 FILLER_165_205 ();
 fill_4 FILLER_165_217 ();
 fill_2 FILLER_165_221 ();
 fill_1 FILLER_165_223 ();
 decap_12 FILLER_165_225 ();
 decap_12 FILLER_165_237 ();
 fill_4 FILLER_165_284 ();
 fill_1 FILLER_165_300 ();
 fill_2 FILLER_165_328 ();
 fill_1 FILLER_165_330 ();
 fill_2 FILLER_165_373 ();
 fill_1 FILLER_165_375 ();
 fill_1 FILLER_165_381 ();
 fill_2 FILLER_165_390 ();
 fill_4 FILLER_165_393 ();
 fill_2 FILLER_165_397 ();
 decap_12 FILLER_165_464 ();
 fill_8 FILLER_165_476 ();
 decap_12 FILLER_165_505 ();
 decap_12 FILLER_165_517 ();
 fill_4 FILLER_165_529 ();
 fill_2 FILLER_165_533 ();
 fill_1 FILLER_165_535 ();
 decap_12 FILLER_165_542 ();
 fill_4 FILLER_165_554 ();
 fill_2 FILLER_165_558 ();
 decap_12 FILLER_165_561 ();
 decap_12 FILLER_165_573 ();
 decap_12 FILLER_165_585 ();
 decap_12 FILLER_165_597 ();
 fill_1 FILLER_165_609 ();
 decap_12 FILLER_165_617 ();
 decap_12 FILLER_165_629 ();
 decap_12 FILLER_165_641 ();
 decap_12 FILLER_165_653 ();
 fill_4 FILLER_165_665 ();
 fill_2 FILLER_165_669 ();
 fill_1 FILLER_165_671 ();
 decap_12 FILLER_165_681 ();
 decap_12 FILLER_165_693 ();
 decap_12 FILLER_165_705 ();
 fill_8 FILLER_165_717 ();
 fill_2 FILLER_165_725 ();
 fill_1 FILLER_165_727 ();
 fill_1 FILLER_165_729 ();
 fill_1 FILLER_165_783 ();
 fill_8 FILLER_165_813 ();
 fill_2 FILLER_165_827 ();
 fill_8 FILLER_165_832 ();
 fill_4 FILLER_165_841 ();
 fill_1 FILLER_165_845 ();
 fill_2 FILLER_165_849 ();
 fill_4 FILLER_165_868 ();
 fill_2 FILLER_165_872 ();
 fill_1 FILLER_165_874 ();
 fill_1 FILLER_165_883 ();
 fill_2 FILLER_165_893 ();
 fill_1 FILLER_165_895 ();
 decap_12 FILLER_165_902 ();
 decap_12 FILLER_165_914 ();
 decap_12 FILLER_165_926 ();
 decap_12 FILLER_165_938 ();
 fill_2 FILLER_165_950 ();
 decap_12 FILLER_165_953 ();
 decap_12 FILLER_165_965 ();
 decap_12 FILLER_165_977 ();
 decap_12 FILLER_165_989 ();
 fill_4 FILLER_165_1001 ();
 fill_2 FILLER_165_1005 ();
 fill_1 FILLER_165_1007 ();
 decap_12 FILLER_165_1009 ();
 decap_12 FILLER_165_1021 ();
 fill_4 FILLER_165_1033 ();
 fill_1 FILLER_165_1037 ();
 decap_12 FILLER_166_5 ();
 fill_8 FILLER_166_17 ();
 fill_2 FILLER_166_25 ();
 fill_1 FILLER_166_27 ();
 decap_12 FILLER_166_29 ();
 decap_12 FILLER_166_41 ();
 decap_12 FILLER_166_53 ();
 decap_12 FILLER_166_65 ();
 fill_4 FILLER_166_77 ();
 fill_2 FILLER_166_81 ();
 fill_1 FILLER_166_83 ();
 decap_12 FILLER_166_85 ();
 decap_12 FILLER_166_97 ();
 decap_12 FILLER_166_109 ();
 decap_12 FILLER_166_121 ();
 fill_4 FILLER_166_133 ();
 fill_2 FILLER_166_137 ();
 fill_1 FILLER_166_139 ();
 decap_12 FILLER_166_141 ();
 decap_12 FILLER_166_153 ();
 decap_12 FILLER_166_165 ();
 decap_12 FILLER_166_177 ();
 fill_4 FILLER_166_189 ();
 fill_2 FILLER_166_193 ();
 fill_1 FILLER_166_195 ();
 decap_12 FILLER_166_197 ();
 decap_12 FILLER_166_209 ();
 decap_12 FILLER_166_221 ();
 decap_12 FILLER_166_233 ();
 fill_4 FILLER_166_245 ();
 fill_2 FILLER_166_249 ();
 fill_1 FILLER_166_251 ();
 fill_2 FILLER_166_253 ();
 fill_4 FILLER_166_309 ();
 fill_2 FILLER_166_313 ();
 fill_2 FILLER_166_320 ();
 fill_4 FILLER_166_330 ();
 fill_4 FILLER_166_415 ();
 fill_1 FILLER_166_419 ();
 fill_1 FILLER_166_467 ();
 fill_4 FILLER_166_477 ();
 fill_1 FILLER_166_481 ();
 decap_12 FILLER_166_514 ();
 fill_4 FILLER_166_526 ();
 fill_2 FILLER_166_530 ();
 decap_12 FILLER_166_533 ();
 fill_4 FILLER_166_545 ();
 fill_2 FILLER_166_549 ();
 fill_1 FILLER_166_551 ();
 decap_12 FILLER_166_555 ();
 decap_12 FILLER_166_573 ();
 fill_2 FILLER_166_585 ();
 fill_1 FILLER_166_587 ();
 fill_1 FILLER_166_589 ();
 decap_12 FILLER_166_596 ();
 decap_12 FILLER_166_608 ();
 decap_12 FILLER_166_620 ();
 decap_12 FILLER_166_632 ();
 fill_4 FILLER_166_650 ();
 decap_12 FILLER_166_678 ();
 fill_8 FILLER_166_690 ();
 fill_2 FILLER_166_698 ();
 decap_12 FILLER_166_701 ();
 decap_12 FILLER_166_713 ();
 decap_12 FILLER_166_725 ();
 fill_4 FILLER_166_737 ();
 fill_1 FILLER_166_741 ();
 fill_4 FILLER_166_745 ();
 fill_1 FILLER_166_749 ();
 fill_2 FILLER_166_754 ();
 fill_4 FILLER_166_757 ();
 fill_2 FILLER_166_780 ();
 fill_2 FILLER_166_802 ();
 fill_4 FILLER_166_807 ();
 fill_1 FILLER_166_811 ();
 fill_2 FILLER_166_813 ();
 fill_1 FILLER_166_815 ();
 fill_8 FILLER_166_860 ();
 fill_4 FILLER_166_886 ();
 decap_12 FILLER_166_901 ();
 fill_8 FILLER_166_913 ();
 fill_2 FILLER_166_921 ();
 fill_1 FILLER_166_923 ();
 decap_12 FILLER_166_925 ();
 decap_12 FILLER_166_937 ();
 decap_12 FILLER_166_949 ();
 decap_12 FILLER_166_961 ();
 fill_4 FILLER_166_973 ();
 fill_2 FILLER_166_977 ();
 fill_1 FILLER_166_979 ();
 decap_12 FILLER_166_981 ();
 decap_12 FILLER_166_993 ();
 decap_12 FILLER_166_1005 ();
 decap_12 FILLER_166_1017 ();
 fill_4 FILLER_166_1029 ();
 fill_2 FILLER_166_1033 ();
 fill_1 FILLER_166_1035 ();
 fill_1 FILLER_166_1037 ();
 decap_12 FILLER_167_5 ();
 decap_12 FILLER_167_17 ();
 decap_12 FILLER_167_29 ();
 decap_12 FILLER_167_41 ();
 fill_2 FILLER_167_53 ();
 fill_1 FILLER_167_55 ();
 decap_12 FILLER_167_57 ();
 decap_12 FILLER_167_69 ();
 decap_12 FILLER_167_81 ();
 decap_12 FILLER_167_93 ();
 fill_4 FILLER_167_105 ();
 fill_2 FILLER_167_109 ();
 fill_1 FILLER_167_111 ();
 decap_12 FILLER_167_113 ();
 decap_12 FILLER_167_125 ();
 decap_12 FILLER_167_137 ();
 decap_12 FILLER_167_149 ();
 fill_4 FILLER_167_161 ();
 fill_2 FILLER_167_165 ();
 fill_1 FILLER_167_167 ();
 decap_12 FILLER_167_169 ();
 decap_12 FILLER_167_181 ();
 decap_12 FILLER_167_193 ();
 decap_12 FILLER_167_205 ();
 fill_4 FILLER_167_217 ();
 fill_2 FILLER_167_221 ();
 fill_1 FILLER_167_223 ();
 decap_12 FILLER_167_225 ();
 decap_12 FILLER_167_237 ();
 fill_8 FILLER_167_249 ();
 fill_2 FILLER_167_257 ();
 decap_12 FILLER_167_264 ();
 fill_4 FILLER_167_276 ();
 fill_2 FILLER_167_281 ();
 decap_12 FILLER_167_290 ();
 fill_4 FILLER_167_332 ();
 fill_2 FILLER_167_346 ();
 fill_4 FILLER_167_380 ();
 fill_4 FILLER_167_393 ();
 fill_2 FILLER_167_397 ();
 fill_1 FILLER_167_408 ();
 fill_4 FILLER_167_441 ();
 fill_2 FILLER_167_445 ();
 fill_1 FILLER_167_447 ();
 fill_8 FILLER_167_449 ();
 fill_1 FILLER_167_477 ();
 fill_1 FILLER_167_486 ();
 decap_12 FILLER_167_490 ();
 fill_2 FILLER_167_502 ();
 fill_4 FILLER_167_505 ();
 fill_2 FILLER_167_509 ();
 fill_1 FILLER_167_511 ();
 decap_12 FILLER_167_515 ();
 fill_2 FILLER_167_527 ();
 fill_1 FILLER_167_529 ();
 decap_12 FILLER_167_535 ();
 fill_4 FILLER_167_547 ();
 fill_2 FILLER_167_557 ();
 fill_1 FILLER_167_559 ();
 fill_4 FILLER_167_561 ();
 fill_2 FILLER_167_565 ();
 decap_12 FILLER_167_573 ();
 decap_12 FILLER_167_585 ();
 decap_12 FILLER_167_597 ();
 fill_4 FILLER_167_609 ();
 fill_2 FILLER_167_613 ();
 fill_1 FILLER_167_615 ();
 decap_12 FILLER_167_617 ();
 fill_2 FILLER_167_629 ();
 fill_4 FILLER_167_634 ();
 fill_2 FILLER_167_638 ();
 fill_1 FILLER_167_640 ();
 fill_8 FILLER_167_664 ();
 decap_12 FILLER_167_673 ();
 decap_12 FILLER_167_685 ();
 decap_12 FILLER_167_697 ();
 decap_12 FILLER_167_709 ();
 fill_4 FILLER_167_721 ();
 fill_2 FILLER_167_725 ();
 fill_1 FILLER_167_727 ();
 decap_12 FILLER_167_729 ();
 fill_4 FILLER_167_741 ();
 fill_1 FILLER_167_745 ();
 fill_8 FILLER_167_774 ();
 fill_2 FILLER_167_782 ();
 fill_1 FILLER_167_785 ();
 fill_8 FILLER_167_789 ();
 fill_2 FILLER_167_797 ();
 fill_1 FILLER_167_799 ();
 fill_4 FILLER_167_819 ();
 fill_2 FILLER_167_823 ();
 fill_2 FILLER_167_834 ();
 fill_1 FILLER_167_836 ();
 fill_2 FILLER_167_841 ();
 fill_4 FILLER_167_879 ();
 fill_1 FILLER_167_883 ();
 fill_2 FILLER_167_894 ();
 decap_12 FILLER_167_897 ();
 decap_12 FILLER_167_909 ();
 decap_12 FILLER_167_921 ();
 decap_12 FILLER_167_933 ();
 fill_4 FILLER_167_945 ();
 fill_2 FILLER_167_949 ();
 fill_1 FILLER_167_951 ();
 decap_12 FILLER_167_953 ();
 decap_12 FILLER_167_965 ();
 decap_12 FILLER_167_977 ();
 decap_12 FILLER_167_989 ();
 fill_4 FILLER_167_1001 ();
 fill_2 FILLER_167_1005 ();
 fill_1 FILLER_167_1007 ();
 decap_12 FILLER_167_1009 ();
 decap_12 FILLER_167_1021 ();
 fill_4 FILLER_167_1033 ();
 fill_1 FILLER_167_1037 ();
 decap_12 FILLER_168_3 ();
 decap_12 FILLER_168_15 ();
 fill_1 FILLER_168_27 ();
 decap_12 FILLER_168_29 ();
 decap_12 FILLER_168_41 ();
 decap_12 FILLER_168_53 ();
 decap_12 FILLER_168_65 ();
 fill_4 FILLER_168_77 ();
 fill_2 FILLER_168_81 ();
 fill_1 FILLER_168_83 ();
 decap_12 FILLER_168_85 ();
 decap_12 FILLER_168_97 ();
 decap_12 FILLER_168_109 ();
 decap_12 FILLER_168_121 ();
 fill_4 FILLER_168_133 ();
 fill_2 FILLER_168_137 ();
 fill_1 FILLER_168_139 ();
 decap_12 FILLER_168_141 ();
 decap_12 FILLER_168_153 ();
 decap_12 FILLER_168_165 ();
 decap_12 FILLER_168_177 ();
 fill_4 FILLER_168_189 ();
 fill_2 FILLER_168_193 ();
 fill_1 FILLER_168_195 ();
 decap_12 FILLER_168_197 ();
 decap_12 FILLER_168_209 ();
 decap_12 FILLER_168_221 ();
 decap_12 FILLER_168_233 ();
 fill_4 FILLER_168_245 ();
 fill_2 FILLER_168_249 ();
 fill_1 FILLER_168_251 ();
 decap_12 FILLER_168_253 ();
 decap_12 FILLER_168_265 ();
 decap_12 FILLER_168_277 ();
 decap_12 FILLER_168_289 ();
 fill_4 FILLER_168_301 ();
 fill_2 FILLER_168_305 ();
 fill_1 FILLER_168_307 ();
 fill_2 FILLER_168_309 ();
 fill_1 FILLER_168_325 ();
 fill_1 FILLER_168_350 ();
 fill_2 FILLER_168_362 ();
 fill_1 FILLER_168_365 ();
 fill_1 FILLER_168_387 ();
 fill_2 FILLER_168_408 ();
 fill_1 FILLER_168_410 ();
 fill_8 FILLER_168_447 ();
 fill_2 FILLER_168_455 ();
 fill_1 FILLER_168_475 ();
 decap_12 FILLER_168_497 ();
 decap_12 FILLER_168_509 ();
 fill_8 FILLER_168_521 ();
 fill_2 FILLER_168_529 ();
 fill_1 FILLER_168_531 ();
 decap_12 FILLER_168_533 ();
 decap_12 FILLER_168_545 ();
 decap_12 FILLER_168_557 ();
 decap_12 FILLER_168_569 ();
 fill_4 FILLER_168_581 ();
 fill_2 FILLER_168_585 ();
 fill_1 FILLER_168_587 ();
 fill_4 FILLER_168_595 ();
 fill_2 FILLER_168_599 ();
 fill_8 FILLER_168_606 ();
 fill_2 FILLER_168_614 ();
 decap_12 FILLER_168_620 ();
 decap_12 FILLER_168_632 ();
 decap_12 FILLER_168_645 ();
 decap_12 FILLER_168_657 ();
 decap_12 FILLER_168_669 ();
 decap_12 FILLER_168_681 ();
 fill_4 FILLER_168_693 ();
 fill_2 FILLER_168_697 ();
 fill_1 FILLER_168_699 ();
 decap_12 FILLER_168_701 ();
 decap_12 FILLER_168_713 ();
 fill_2 FILLER_168_725 ();
 fill_8 FILLER_168_748 ();
 decap_12 FILLER_168_757 ();
 fill_1 FILLER_168_769 ();
 fill_1 FILLER_168_791 ();
 fill_1 FILLER_168_813 ();
 decap_12 FILLER_168_894 ();
 decap_12 FILLER_168_906 ();
 fill_4 FILLER_168_918 ();
 fill_2 FILLER_168_922 ();
 decap_12 FILLER_168_925 ();
 decap_12 FILLER_168_937 ();
 decap_12 FILLER_168_949 ();
 decap_12 FILLER_168_961 ();
 fill_4 FILLER_168_973 ();
 fill_2 FILLER_168_977 ();
 fill_1 FILLER_168_979 ();
 decap_12 FILLER_168_981 ();
 decap_12 FILLER_168_993 ();
 decap_12 FILLER_168_1005 ();
 decap_12 FILLER_168_1017 ();
 fill_4 FILLER_168_1029 ();
 fill_2 FILLER_168_1033 ();
 fill_1 FILLER_168_1035 ();
 fill_1 FILLER_168_1037 ();
 decap_12 FILLER_169_3 ();
 decap_12 FILLER_169_15 ();
 decap_12 FILLER_169_27 ();
 decap_12 FILLER_169_39 ();
 fill_4 FILLER_169_51 ();
 fill_1 FILLER_169_55 ();
 decap_12 FILLER_169_57 ();
 decap_12 FILLER_169_69 ();
 decap_12 FILLER_169_81 ();
 decap_12 FILLER_169_93 ();
 fill_4 FILLER_169_105 ();
 fill_2 FILLER_169_109 ();
 fill_1 FILLER_169_111 ();
 decap_12 FILLER_169_113 ();
 decap_12 FILLER_169_125 ();
 decap_12 FILLER_169_137 ();
 decap_12 FILLER_169_149 ();
 fill_4 FILLER_169_161 ();
 fill_2 FILLER_169_165 ();
 fill_1 FILLER_169_167 ();
 decap_12 FILLER_169_169 ();
 decap_12 FILLER_169_181 ();
 decap_12 FILLER_169_193 ();
 decap_12 FILLER_169_205 ();
 fill_4 FILLER_169_217 ();
 fill_2 FILLER_169_221 ();
 fill_1 FILLER_169_223 ();
 decap_12 FILLER_169_225 ();
 decap_12 FILLER_169_237 ();
 decap_12 FILLER_169_249 ();
 decap_12 FILLER_169_261 ();
 fill_4 FILLER_169_273 ();
 fill_2 FILLER_169_277 ();
 fill_1 FILLER_169_279 ();
 decap_12 FILLER_169_281 ();
 decap_12 FILLER_169_293 ();
 fill_2 FILLER_169_305 ();
 fill_2 FILLER_169_328 ();
 fill_1 FILLER_169_330 ();
 fill_2 FILLER_169_346 ();
 fill_2 FILLER_169_369 ();
 fill_4 FILLER_169_393 ();
 fill_2 FILLER_169_397 ();
 fill_2 FILLER_169_456 ();
 fill_4 FILLER_169_497 ();
 fill_2 FILLER_169_501 ();
 fill_1 FILLER_169_503 ();
 decap_12 FILLER_169_513 ();
 decap_12 FILLER_169_525 ();
 decap_12 FILLER_169_537 ();
 fill_4 FILLER_169_549 ();
 fill_1 FILLER_169_553 ();
 fill_2 FILLER_169_557 ();
 fill_1 FILLER_169_559 ();
 decap_12 FILLER_169_561 ();
 decap_12 FILLER_169_573 ();
 decap_12 FILLER_169_585 ();
 decap_12 FILLER_169_597 ();
 fill_4 FILLER_169_609 ();
 fill_2 FILLER_169_613 ();
 fill_1 FILLER_169_615 ();
 decap_12 FILLER_169_617 ();
 decap_12 FILLER_169_629 ();
 fill_2 FILLER_169_649 ();
 fill_1 FILLER_169_659 ();
 fill_4 FILLER_169_668 ();
 fill_1 FILLER_169_697 ();
 fill_1 FILLER_169_706 ();
 decap_12 FILLER_169_715 ();
 fill_1 FILLER_169_727 ();
 fill_2 FILLER_169_729 ();
 fill_4 FILLER_169_734 ();
 fill_2 FILLER_169_738 ();
 fill_1 FILLER_169_740 ();
 decap_12 FILLER_169_757 ();
 decap_12 FILLER_169_769 ();
 fill_2 FILLER_169_781 ();
 fill_1 FILLER_169_783 ();
 fill_1 FILLER_169_788 ();
 fill_1 FILLER_169_810 ();
 decap_12 FILLER_169_815 ();
 fill_4 FILLER_169_827 ();
 fill_4 FILLER_169_835 ();
 fill_1 FILLER_169_839 ();
 fill_4 FILLER_169_891 ();
 fill_1 FILLER_169_895 ();
 decap_12 FILLER_169_897 ();
 decap_12 FILLER_169_909 ();
 decap_12 FILLER_169_921 ();
 decap_12 FILLER_169_933 ();
 fill_4 FILLER_169_945 ();
 fill_2 FILLER_169_949 ();
 fill_1 FILLER_169_951 ();
 decap_12 FILLER_169_953 ();
 decap_12 FILLER_169_965 ();
 decap_12 FILLER_169_977 ();
 decap_12 FILLER_169_989 ();
 fill_4 FILLER_169_1001 ();
 fill_2 FILLER_169_1005 ();
 fill_1 FILLER_169_1007 ();
 decap_12 FILLER_169_1009 ();
 decap_12 FILLER_169_1021 ();
 fill_4 FILLER_169_1033 ();
 fill_1 FILLER_169_1037 ();
 decap_12 FILLER_170_3 ();
 decap_12 FILLER_170_15 ();
 fill_1 FILLER_170_27 ();
 decap_12 FILLER_170_29 ();
 decap_12 FILLER_170_41 ();
 decap_12 FILLER_170_53 ();
 decap_12 FILLER_170_65 ();
 fill_4 FILLER_170_77 ();
 fill_2 FILLER_170_81 ();
 fill_1 FILLER_170_83 ();
 decap_12 FILLER_170_85 ();
 decap_12 FILLER_170_97 ();
 decap_12 FILLER_170_109 ();
 decap_12 FILLER_170_121 ();
 fill_4 FILLER_170_133 ();
 fill_2 FILLER_170_137 ();
 fill_1 FILLER_170_139 ();
 decap_12 FILLER_170_141 ();
 decap_12 FILLER_170_153 ();
 decap_12 FILLER_170_165 ();
 decap_12 FILLER_170_177 ();
 fill_4 FILLER_170_189 ();
 fill_2 FILLER_170_193 ();
 fill_1 FILLER_170_195 ();
 decap_12 FILLER_170_197 ();
 decap_12 FILLER_170_209 ();
 decap_12 FILLER_170_221 ();
 decap_12 FILLER_170_233 ();
 fill_4 FILLER_170_245 ();
 fill_2 FILLER_170_249 ();
 fill_1 FILLER_170_251 ();
 decap_12 FILLER_170_253 ();
 decap_12 FILLER_170_265 ();
 decap_12 FILLER_170_277 ();
 decap_12 FILLER_170_289 ();
 fill_4 FILLER_170_301 ();
 fill_2 FILLER_170_305 ();
 fill_1 FILLER_170_307 ();
 fill_2 FILLER_170_309 ();
 fill_2 FILLER_170_337 ();
 fill_1 FILLER_170_363 ();
 fill_2 FILLER_170_365 ();
 fill_1 FILLER_170_367 ();
 fill_4 FILLER_170_377 ();
 fill_2 FILLER_170_417 ();
 fill_1 FILLER_170_419 ();
 fill_2 FILLER_170_430 ();
 fill_1 FILLER_170_432 ();
 fill_1 FILLER_170_453 ();
 decap_12 FILLER_170_497 ();
 fill_8 FILLER_170_509 ();
 fill_2 FILLER_170_517 ();
 fill_1 FILLER_170_519 ();
 fill_4 FILLER_170_526 ();
 fill_2 FILLER_170_530 ();
 fill_8 FILLER_170_533 ();
 decap_12 FILLER_170_547 ();
 fill_8 FILLER_170_559 ();
 fill_1 FILLER_170_567 ();
 fill_8 FILLER_170_579 ();
 fill_1 FILLER_170_587 ();
 decap_12 FILLER_170_589 ();
 fill_8 FILLER_170_601 ();
 fill_2 FILLER_170_617 ();
 fill_2 FILLER_170_627 ();
 fill_4 FILLER_170_637 ();
 fill_2 FILLER_170_641 ();
 fill_1 FILLER_170_643 ();
 decap_12 FILLER_170_645 ();
 decap_12 FILLER_170_657 ();
 decap_12 FILLER_170_669 ();
 decap_12 FILLER_170_681 ();
 fill_4 FILLER_170_693 ();
 fill_2 FILLER_170_697 ();
 fill_1 FILLER_170_699 ();
 decap_12 FILLER_170_701 ();
 decap_12 FILLER_170_713 ();
 decap_12 FILLER_170_725 ();
 decap_12 FILLER_170_737 ();
 fill_4 FILLER_170_749 ();
 fill_2 FILLER_170_753 ();
 fill_1 FILLER_170_755 ();
 decap_12 FILLER_170_757 ();
 decap_12 FILLER_170_769 ();
 decap_12 FILLER_170_781 ();
 fill_8 FILLER_170_793 ();
 fill_2 FILLER_170_801 ();
 fill_4 FILLER_170_806 ();
 fill_2 FILLER_170_810 ();
 decap_12 FILLER_170_813 ();
 decap_12 FILLER_170_825 ();
 fill_2 FILLER_170_837 ();
 fill_1 FILLER_170_839 ();
 decap_12 FILLER_170_893 ();
 decap_12 FILLER_170_905 ();
 fill_4 FILLER_170_917 ();
 fill_2 FILLER_170_921 ();
 fill_1 FILLER_170_923 ();
 decap_12 FILLER_170_925 ();
 decap_12 FILLER_170_937 ();
 decap_12 FILLER_170_949 ();
 decap_12 FILLER_170_961 ();
 fill_4 FILLER_170_973 ();
 fill_2 FILLER_170_977 ();
 fill_1 FILLER_170_979 ();
 decap_12 FILLER_170_981 ();
 decap_12 FILLER_170_993 ();
 decap_12 FILLER_170_1005 ();
 decap_12 FILLER_170_1017 ();
 fill_2 FILLER_170_1029 ();
 fill_1 FILLER_170_1031 ();
 fill_2 FILLER_170_1034 ();
 fill_1 FILLER_170_1037 ();
 decap_12 FILLER_171_3 ();
 decap_12 FILLER_171_15 ();
 fill_1 FILLER_171_27 ();
 decap_12 FILLER_171_29 ();
 decap_12 FILLER_171_41 ();
 fill_2 FILLER_171_53 ();
 fill_1 FILLER_171_55 ();
 decap_12 FILLER_171_57 ();
 decap_12 FILLER_171_69 ();
 fill_2 FILLER_171_81 ();
 fill_1 FILLER_171_83 ();
 decap_12 FILLER_171_85 ();
 decap_12 FILLER_171_97 ();
 fill_2 FILLER_171_109 ();
 fill_1 FILLER_171_111 ();
 decap_12 FILLER_171_113 ();
 decap_12 FILLER_171_125 ();
 fill_2 FILLER_171_137 ();
 fill_1 FILLER_171_139 ();
 decap_12 FILLER_171_141 ();
 decap_12 FILLER_171_153 ();
 fill_2 FILLER_171_165 ();
 fill_1 FILLER_171_167 ();
 decap_12 FILLER_171_169 ();
 decap_12 FILLER_171_181 ();
 fill_2 FILLER_171_193 ();
 fill_1 FILLER_171_195 ();
 decap_12 FILLER_171_197 ();
 decap_12 FILLER_171_209 ();
 fill_2 FILLER_171_221 ();
 fill_1 FILLER_171_223 ();
 decap_12 FILLER_171_225 ();
 decap_12 FILLER_171_237 ();
 fill_2 FILLER_171_249 ();
 fill_1 FILLER_171_251 ();
 decap_12 FILLER_171_253 ();
 decap_12 FILLER_171_265 ();
 fill_2 FILLER_171_277 ();
 fill_1 FILLER_171_279 ();
 decap_12 FILLER_171_281 ();
 decap_12 FILLER_171_293 ();
 fill_2 FILLER_171_305 ();
 fill_1 FILLER_171_307 ();
 decap_12 FILLER_171_309 ();
 fill_1 FILLER_171_321 ();
 fill_8 FILLER_171_337 ();
 fill_2 FILLER_171_350 ();
 fill_2 FILLER_171_361 ();
 fill_1 FILLER_171_363 ();
 fill_1 FILLER_171_391 ();
 fill_2 FILLER_171_393 ();
 fill_1 FILLER_171_395 ();
 fill_4 FILLER_171_421 ();
 fill_2 FILLER_171_425 ();
 fill_2 FILLER_171_445 ();
 fill_1 FILLER_171_447 ();
 fill_4 FILLER_171_449 ();
 fill_1 FILLER_171_453 ();
 fill_8 FILLER_171_460 ();
 fill_1 FILLER_171_468 ();
 fill_2 FILLER_171_474 ();
 decap_12 FILLER_171_477 ();
 fill_4 FILLER_171_489 ();
 fill_2 FILLER_171_493 ();
 fill_1 FILLER_171_495 ();
 decap_12 FILLER_171_513 ();
 fill_4 FILLER_171_525 ();
 fill_2 FILLER_171_529 ();
 fill_1 FILLER_171_531 ();
 decap_12 FILLER_171_533 ();
 fill_4 FILLER_171_545 ();
 fill_1 FILLER_171_549 ();
 fill_2 FILLER_171_558 ();
 decap_12 FILLER_171_561 ();
 decap_12 FILLER_171_573 ();
 fill_2 FILLER_171_585 ();
 fill_1 FILLER_171_587 ();
 fill_2 FILLER_171_597 ();
 fill_8 FILLER_171_607 ();
 fill_1 FILLER_171_615 ();
 decap_12 FILLER_171_617 ();
 decap_12 FILLER_171_629 ();
 fill_2 FILLER_171_641 ();
 fill_1 FILLER_171_643 ();
 decap_12 FILLER_171_645 ();
 decap_12 FILLER_171_657 ();
 fill_2 FILLER_171_669 ();
 fill_1 FILLER_171_671 ();
 decap_12 FILLER_171_673 ();
 decap_12 FILLER_171_685 ();
 fill_2 FILLER_171_697 ();
 fill_1 FILLER_171_699 ();
 decap_12 FILLER_171_701 ();
 decap_12 FILLER_171_713 ();
 fill_2 FILLER_171_725 ();
 fill_1 FILLER_171_727 ();
 decap_12 FILLER_171_729 ();
 decap_12 FILLER_171_741 ();
 fill_2 FILLER_171_753 ();
 fill_1 FILLER_171_755 ();
 decap_12 FILLER_171_757 ();
 decap_12 FILLER_171_769 ();
 fill_2 FILLER_171_781 ();
 fill_1 FILLER_171_783 ();
 decap_12 FILLER_171_785 ();
 decap_12 FILLER_171_797 ();
 fill_2 FILLER_171_809 ();
 fill_1 FILLER_171_811 ();
 decap_12 FILLER_171_813 ();
 decap_12 FILLER_171_825 ();
 fill_2 FILLER_171_837 ();
 fill_1 FILLER_171_839 ();
 decap_12 FILLER_171_841 ();
 fill_4 FILLER_171_853 ();
 fill_2 FILLER_171_861 ();
 fill_2 FILLER_171_866 ();
 fill_8 FILLER_171_888 ();
 decap_12 FILLER_171_897 ();
 decap_12 FILLER_171_909 ();
 fill_2 FILLER_171_921 ();
 fill_1 FILLER_171_923 ();
 decap_12 FILLER_171_925 ();
 decap_12 FILLER_171_937 ();
 fill_2 FILLER_171_949 ();
 fill_1 FILLER_171_951 ();
 decap_12 FILLER_171_953 ();
 decap_12 FILLER_171_965 ();
 fill_2 FILLER_171_977 ();
 fill_1 FILLER_171_979 ();
 decap_12 FILLER_171_981 ();
 decap_12 FILLER_171_993 ();
 fill_2 FILLER_171_1005 ();
 fill_1 FILLER_171_1007 ();
 decap_12 FILLER_171_1009 ();
 fill_1 FILLER_171_1021 ();
 fill_1 FILLER_171_1037 ();

endmodule
